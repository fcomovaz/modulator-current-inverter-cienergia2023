LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY Ratio1 IS
    PORT (
        clk : IN STD_LOGIC;
        rst : IN STD_LOGIC;
        adc_cum_sum : IN UNSIGNED(23 DOWNTO 0);
        lut_value : OUT INTEGER RANGE 0 TO 18000
    );
END ENTITY Ratio1;

ARCHITECTURE main OF Ratio1 IS
    -- LUT definition with 11 elements (index 0 to 10)
    TYPE LUT_TYPE IS ARRAY (0 TO 71999) OF INTEGER RANGE 0 TO 72000;
    CONSTANT lut_values : LUT_TYPE := (36000, 35978, 35978, 35978, 35951, 35951, 35951, 35929, 35929, 35929, 35902, 35902, 35880, 35880, 35880, 35853, 35853, 35853, 35831, 35831, 35831, 35804, 35804, 35804, 35782, 35782, 35782, 35755, 35755, 35755, 35733, 35733, 35706, 35706, 35706, 35684, 35684, 35684, 35657, 35657, 35657, 35635, 35635, 35635, 35608, 35608, 35608, 35586, 35586, 35586, 35559, 35559, 35537, 35537, 35537, 35510, 35510, 35510, 35488, 35488, 35488, 35461, 35461, 35461, 35440, 35440, 35440, 35412, 35412, 35412, 35391, 35391, 35363, 35363, 35363, 35342, 35342, 35342, 35314, 35314, 35314, 35293, 35293, 35293, 35265, 35265, 35265, 35244, 35244, 35244, 35216, 35216, 35195, 35195, 35195, 35167, 35167, 35167, 35146, 35146, 35146, 35118, 35118, 35118, 35097, 35097, 35097, 35069, 35069, 35069, 35048, 35048, 35020, 35020, 35020, 34999, 34999, 34999, 34971, 34971, 34971, 34950, 34950, 34950, 34922, 34922, 34922, 34901, 34901, 34901, 34879, 34879, 34852, 34852, 34852, 34830, 34830, 34830, 34803, 34803, 34803, 34781, 34781, 34781, 34754, 34754, 34754, 34732, 34732, 34732, 34705, 34705, 34683, 34683, 34683, 34656, 34656, 34656, 34634, 34634, 34634, 34607, 34607, 34607, 34585, 34585, 34585, 34558, 34558, 34558, 34536, 34536, 34509, 34509, 34509, 34487, 34487, 34487, 34460, 34460, 34460, 34438, 34438, 34438, 34411, 34411, 34411, 34389, 34389, 34389, 34362, 34362, 34340, 34340, 34340, 34313, 34313, 34313, 34291, 34291, 34291, 34264, 34264, 34264, 34242, 34242, 34242, 34215, 34215, 34215, 34193, 34193, 34166, 34166, 34166, 34144, 34144, 34144, 34117, 34117, 34117, 34095, 34095, 34095, 34068, 34068, 34068, 34046, 34046, 34046, 34019, 34019, 33997, 33997, 33997, 33970, 33970, 33970, 33948, 33948, 33948, 33921, 33921, 33921, 33899, 33899, 33899, 33872, 33872, 33872, 33850, 33850, 33823, 33823, 33823, 33801, 33801, 33801, 33779, 33779, 33779, 33752, 33752, 33752, 33730, 33730, 33730, 33703, 33703, 33703, 33681, 33681, 33654, 33654, 33654, 33632, 33632, 33632, 33605, 33605, 33605, 33583, 33583, 33583, 33556, 33556, 33556, 33534, 33534, 33534, 33507, 33507, 33485, 33485, 33485, 33457, 33457, 33457, 33436, 33436, 33436, 33408, 33408, 33408, 33387, 33387, 33387, 33359, 33359, 33359, 33338, 33338, 33310, 33310, 33310, 33288, 33288, 33288, 33261, 33261, 33261, 33239, 33239, 33239, 33212, 33212, 33212, 33190, 33190, 33190, 33163, 33163, 33141, 33141, 33141, 33114, 33114, 33114, 33092, 33092, 33092, 33065, 33065, 33065, 33043, 33043, 33043, 33016, 33016, 33016, 32994, 32994, 32967, 32967, 32967, 32945, 32945, 32945, 32918, 32918, 32918, 32896, 32896, 32896, 32869, 32869, 32869, 32847, 32847, 32847, 32819, 32819, 32798, 32798, 32798, 32770, 32770, 32770, 32749, 32749, 32749, 32727, 32727, 32727, 32699, 32699, 32699, 32678, 32678, 32678, 32650, 32650, 32650, 32628, 32628, 32601, 32601, 32601, 32579, 32579, 32579, 32552, 32552, 32552, 32530, 32530, 32530, 32503, 32503, 32503, 32481, 32481, 32481, 32454, 32454, 32432, 32432, 32432, 32405, 32405, 32405, 32383, 32383, 32383, 32356, 32356, 32356, 32334, 32334, 32334, 32306, 32306, 32306, 32285, 32285, 32257, 32257, 32257, 32235, 32235, 32235, 32208, 32208, 32208, 32186, 32186, 32186, 32159, 32159, 32159, 32137, 32137, 32137, 32110, 32110, 32088, 32088, 32088, 32061, 32061, 32061, 32039, 32039, 32039, 32011, 32011, 32011, 31990, 31990, 31990, 31962, 31962, 31962, 31940, 31940, 31913, 31913, 31913, 31891, 31891, 31891, 31864, 31864, 31864, 31842, 31842, 31842, 31815, 31815, 31815, 31793, 31793, 31793, 31766, 31766, 31744, 31744, 31744, 31716, 31716, 31716, 31694, 31694, 31694, 31667, 31667, 31667, 31645, 31645, 31645, 31623, 31623, 31623, 31596, 31596, 31574, 31574, 31574, 31547, 31547, 31547, 31525, 31525, 31525, 31498, 31498, 31498, 31476, 31476, 31476, 31448, 31448, 31448, 31426, 31426, 31426, 31399, 31399, 31377, 31377, 31377, 31350, 31350, 31350, 31328, 31328, 31328, 31301, 31301, 31301, 31279, 31279, 31279, 31251, 31251, 31251, 31230, 31230, 31202, 31202, 31202, 31180, 31180, 31180, 31153, 31153, 31153, 31131, 31131, 31131, 31104, 31104, 31104, 31082, 31082, 31082, 31054, 31054, 31032, 31032, 31032, 31005, 31005, 31005, 30983, 30983, 30983, 30956, 30956, 30956, 30934, 30934, 30934, 30906, 30906, 30906, 30885, 30885, 30857, 30857, 30857, 30835, 30835, 30835, 30808, 30808, 30808, 30786, 30786, 30786, 30759, 30759, 30759, 30737, 30737, 30737, 30709, 30709, 30687, 30687, 30687, 30660, 30660, 30660, 30638, 30638, 30638, 30611, 30611, 30611, 30589, 30589, 30589, 30561, 30561, 30561, 30539, 30539, 30539, 30517, 30517, 30490, 30490, 30490, 30468, 30468, 30468, 30441, 30441, 30441, 30419, 30419, 30419, 30391, 30391, 30391, 30369, 30369, 30369, 30342, 30342, 30320, 30320, 30320, 30292, 30292, 30292, 30270, 30270, 30270, 30243, 30243, 30243, 30221, 30221, 30221, 30194, 30194, 30194, 30172, 30172, 30144, 30144, 30144, 30122, 30122, 30122, 30095, 30095, 30095, 30073, 30073, 30073, 30045, 30045, 30045, 30023, 30023, 30023, 29996, 29996, 29974, 29974, 29974, 29947, 29947, 29947, 29925, 29925, 29925, 29897, 29897, 29897, 29875, 29875, 29875, 29848, 29848, 29848, 29826, 29826, 29826, 29798, 29798, 29776, 29776, 29776, 29749, 29749, 29749, 29727, 29727, 29727, 29699, 29699, 29699, 29677, 29677, 29677, 29650, 29650, 29650, 29628, 29628, 29600, 29600, 29600, 29578, 29578, 29578, 29551, 29551, 29551, 29529, 29529, 29529, 29501, 29501, 29501, 29479, 29479, 29479, 29452, 29452, 29430, 29430, 29430, 29408, 29408, 29408, 29380, 29380, 29380, 29358, 29358, 29358, 29331, 29331, 29331, 29309, 29309, 29309, 29281, 29281, 29281, 29259, 29259, 29232, 29232, 29232, 29210, 29210, 29210, 29182, 29182, 29182, 29160, 29160, 29160, 29133, 29133, 29133, 29111, 29111, 29111, 29083, 29083, 29061, 29061, 29061, 29033, 29033, 29033, 29011, 29011, 29011, 28984, 28984, 28984, 28962, 28962, 28962, 28934, 28934, 28934, 28912, 28912, 28912, 28885, 28885, 28863, 28863, 28863, 28835, 28835, 28835, 28813, 28813, 28813, 28785, 28785, 28785, 28763, 28763, 28763, 28736, 28736, 28736, 28714, 28714, 28686, 28686, 28686, 28664, 28664, 28664, 28636, 28636, 28636, 28614, 28614, 28614, 28587, 28587, 28587, 28565, 28565, 28565, 28537, 28537, 28515, 28515, 28515, 28487, 28487, 28487, 28465, 28465, 28465, 28438, 28438, 28438, 28416, 28416, 28416, 28388, 28388, 28388, 28366, 28366, 28366, 28344, 28344, 28316, 28316, 28316, 28294, 28294, 28294, 28267, 28267, 28267, 28244, 28244, 28244, 28217, 28217, 28217, 28195, 28195, 28195, 28167, 28167, 28145, 28145, 28145, 28117, 28117, 28117, 28095, 28095, 28095, 28068, 28068, 28068, 28045, 28045, 28045, 28018, 28018, 28018, 27996, 27996, 27996, 27968, 27968, 27946, 27946, 27946, 27918, 27918, 27918, 27896, 27896, 27896, 27868, 27868, 27868, 27846, 27846, 27846, 27819, 27819, 27819, 27796, 27796, 27769, 27769, 27769, 27747, 27747, 27747, 27719, 27719, 27719, 27697, 27697, 27697, 27669, 27669, 27669, 27647, 27647, 27647, 27619, 27619, 27619, 27597, 27597, 27569, 27569, 27569, 27547, 27547, 27547, 27520, 27520, 27520, 27497, 27497, 27497, 27470, 27470, 27470, 27448, 27448, 27448, 27420, 27420, 27420, 27398, 27398, 27370, 27370, 27370, 27348, 27348, 27348, 27320, 27320, 27320, 27298, 27298, 27298, 27270, 27270, 27270, 27248, 27248, 27248, 27226, 27226, 27198, 27198, 27198, 27176, 27176, 27176, 27148, 27148, 27148, 27126, 27126, 27126, 27098, 27098, 27098, 27076, 27076, 27076, 27048, 27048, 27048, 27026, 27026, 26998, 26998, 26998, 26976, 26976, 26976, 26948, 26948, 26948, 26926, 26926, 26926, 26898, 26898, 26898, 26876, 26876, 26876, 26848, 26848, 26848, 26826, 26826, 26798, 26798, 26798, 26776, 26776, 26776, 26748, 26748, 26748, 26726, 26726, 26726, 26698, 26698, 26698, 26676, 26676, 26676, 26648, 26648, 26626, 26626, 26626, 26598, 26598, 26598, 26575, 26575, 26575, 26548, 26548, 26548, 26525, 26525, 26525, 26498, 26498, 26498, 26475, 26475, 26475, 26447, 26447, 26425, 26425, 26425, 26397, 26397, 26397, 26375, 26375, 26375, 26347, 26347, 26347, 26325, 26325, 26325, 26297, 26297, 26297, 26275, 26275, 26275, 26247, 26247, 26225, 26225, 26225, 26197, 26197, 26197, 26174, 26174, 26174, 26146, 26146, 26146, 26124, 26124, 26124, 26102, 26102, 26102, 26074, 26074, 26074, 26052, 26052, 26024, 26024, 26024, 26001, 26001, 26001, 25973, 25973, 25973, 25951, 25951, 25951, 25923, 25923, 25923, 25901, 25901, 25901, 25873, 25873, 25851, 25851, 25851, 25823, 25823, 25823, 25800, 25800, 25800, 25772, 25772, 25772, 25750, 25750, 25750, 25722, 25722, 25722, 25700, 25700, 25700, 25672, 25672, 25649, 25649, 25649, 25621, 25621, 25621, 25599, 25599, 25599, 25571, 25571, 25571, 25549, 25549, 25549, 25521, 25521, 25521, 25498, 25498, 25498, 25470, 25470, 25448, 25448, 25448, 25420, 25420, 25420, 25398, 25398, 25398, 25370, 25370, 25370, 25347, 25347, 25347, 25319, 25319, 25319, 25297, 25297, 25297, 25269, 25269, 25246, 25246, 25246, 25218, 25218, 25218, 25196, 25196, 25196, 25168, 25168, 25168, 25146, 25146, 25146, 25118, 25118, 25118, 25095, 25095, 25095, 25067, 25067, 25045, 25045, 25045, 25017, 25017, 25017, 24994, 24994, 24994, 24972, 24972, 24972, 24944, 24944, 24944, 24921, 24921, 24921, 24893, 24893, 24893, 24871, 24871, 24843, 24843, 24843, 24820, 24820, 24820, 24792, 24792, 24792, 24770, 24770, 24770, 24741, 24741, 24741, 24719, 24719, 24719, 24691, 24691, 24691, 24668, 24668, 24640, 24640, 24640, 24618, 24618, 24618, 24590, 24590, 24590, 24567, 24567, 24567, 24539, 24539, 24539, 24517, 24517, 24517, 24488, 24488, 24488, 24466, 24466, 24438, 24438, 24438, 24415, 24415, 24415, 24387, 24387, 24387, 24365, 24365, 24365, 24336, 24336, 24336, 24314, 24314, 24314, 24286, 24286, 24286, 24263, 24263, 24263, 24235, 24235, 24212, 24212, 24212, 24184, 24184, 24184, 24162, 24162, 24162, 24134, 24134, 24134, 24111, 24111, 24111, 24083, 24083, 24083, 24060, 24060, 24060, 24032, 24032, 24009, 24009, 24009, 23981, 23981, 23981, 23959, 23959, 23959, 23930, 23930, 23930, 23908, 23908, 23908, 23880, 23880, 23880, 23857, 23857, 23857, 23834, 23834, 23806, 23806, 23806, 23784, 23784, 23784, 23755, 23755, 23755, 23733, 23733, 23733, 23704, 23704, 23704, 23682, 23682, 23682, 23654, 23654, 23654, 23631, 23631, 23603, 23603, 23603, 23580, 23580, 23580, 23552, 23552, 23552, 23529, 23529, 23529, 23501, 23501, 23501, 23478, 23478, 23478, 23450, 23450, 23450, 23427, 23427, 23427, 23399, 23399, 23376, 23376, 23376, 23348, 23348, 23348, 23325, 23325, 23325, 23297, 23297, 23297, 23274, 23274, 23274, 23246, 23246, 23246, 23223, 23223, 23223, 23195, 23195, 23172, 23172, 23172, 23144, 23144, 23144, 23121, 23121, 23121, 23093, 23093, 23093, 23070, 23070, 23070, 23042, 23042, 23042, 23019, 23019, 23019, 22991, 22991, 22991, 22968, 22968, 22940, 22940, 22940, 22917, 22917, 22917, 22888, 22888, 22888, 22866, 22866, 22866, 22837, 22837, 22837, 22815, 22815, 22815, 22786, 22786, 22786, 22763, 22763, 22741, 22741, 22741, 22712, 22712, 22712, 22689, 22689, 22689, 22661, 22661, 22661, 22638, 22638, 22638, 22610, 22610, 22610, 22587, 22587, 22587, 22558, 22558, 22558, 22536, 22536, 22507, 22507, 22507, 22484, 22484, 22484, 22456, 22456, 22456, 22433, 22433, 22433, 22405, 22405, 22405, 22382, 22382, 22382, 22353, 22353, 22353, 22331, 22331, 22331, 22302, 22302, 22279, 22279, 22279, 22251, 22251, 22251, 22228, 22228, 22228, 22199, 22199, 22199, 22176, 22176, 22176, 22148, 22148, 22148, 22125, 22125, 22125, 22097, 22097, 22074, 22074, 22074, 22045, 22045, 22045, 22022, 22022, 22022, 21994, 21994, 21994, 21971, 21971, 21971, 21942, 21942, 21942, 21919, 21919, 21919, 21891, 21891, 21891, 21868, 21868, 21839, 21839, 21839, 21816, 21816, 21816, 21788, 21788, 21788, 21765, 21765, 21765, 21736, 21736, 21736, 21713, 21713, 21713, 21685, 21685, 21685, 21662, 21662, 21662, 21633, 21633, 21610, 21610, 21610, 21587, 21587, 21587, 21559, 21559, 21559, 21536, 21536, 21536, 21507, 21507, 21507, 21484, 21484, 21484, 21455, 21455, 21455, 21432, 21432, 21432, 21404, 21404, 21381, 21381, 21381, 21352, 21352, 21352, 21329, 21329, 21329, 21300, 21300, 21300, 21277, 21277, 21277, 21249, 21249, 21249, 21226, 21226, 21226, 21197, 21197, 21197, 21174, 21174, 21145, 21145, 21145, 21122, 21122, 21122, 21093, 21093, 21093, 21070, 21070, 21070, 21042, 21042, 21042, 21019, 21019, 21019, 20990, 20990, 20990, 20967, 20967, 20967, 20938, 20938, 20915, 20915, 20915, 20886, 20886, 20886, 20863, 20863, 20863, 20834, 20834, 20834, 20811, 20811, 20811, 20782, 20782, 20782, 20759, 20759, 20759, 20731, 20731, 20731, 20708, 20708, 20679, 20679, 20679, 20656, 20656, 20656, 20627, 20627, 20627, 20604, 20604, 20604, 20575, 20575, 20575, 20552, 20552, 20552, 20523, 20523, 20523, 20500, 20500, 20500, 20471, 20471, 20471, 20448, 20448, 20425, 20425, 20425, 20396, 20396, 20396, 20373, 20373, 20373, 20344, 20344, 20344, 20320, 20320, 20320, 20292, 20292, 20292, 20268, 20268, 20268, 20239, 20239, 20239, 20216, 20216, 20187, 20187, 20187, 20164, 20164, 20164, 20135, 20135, 20135, 20112, 20112, 20112, 20083, 20083, 20083, 20060, 20060, 20060, 20031, 20031, 20031, 20008, 20008, 20008, 19979, 19979, 19955, 19955, 19955, 19926, 19926, 19926, 19903, 19903, 19903, 19874, 19874, 19874, 19851, 19851, 19851, 19822, 19822, 19822, 19799, 19799, 19799, 19770, 19770, 19770, 19746, 19746, 19746, 19717, 19717, 19694, 19694, 19694, 19665, 19665, 19665, 19642, 19642, 19642, 19613, 19613, 19613, 19589, 19589, 19589, 19560, 19560, 19560, 19537, 19537, 19537, 19508, 19508, 19508, 19485, 19485, 19485, 19456, 19456, 19432, 19432, 19432, 19403, 19403, 19403, 19380, 19380, 19380, 19351, 19351, 19351, 19327, 19327, 19327, 19298, 19298, 19298, 19275, 19275, 19275, 19252, 19252, 19252, 19222, 19222, 19199, 19199, 19199, 19170, 19170, 19170, 19146, 19146, 19146, 19117, 19117, 19117, 19094, 19094, 19094, 19065, 19065, 19065, 19041, 19041, 19041, 19012, 19012, 19012, 18989, 18989, 18989, 18959, 18959, 18936, 18936, 18936, 18907, 18907, 18907, 18883, 18883, 18883, 18854, 18854, 18854, 18831, 18831, 18831, 18801, 18801, 18801, 18778, 18778, 18778, 18749, 18749, 18749, 18725, 18725, 18725, 18696, 18696, 18673, 18673, 18673, 18643, 18643, 18643, 18620, 18620, 18620, 18590, 18590, 18590, 18567, 18567, 18567, 18538, 18538, 18538, 18514, 18514, 18514, 18485, 18485, 18485, 18461, 18461, 18461, 18432, 18432, 18432, 18409, 18409, 18379, 18379, 18379, 18356, 18356, 18356, 18326, 18326, 18326, 18303, 18303, 18303, 18273, 18273, 18273, 18250, 18250, 18250, 18220, 18220, 18220, 18197, 18197, 18197, 18167, 18167, 18167, 18144, 18144, 18120, 18120, 18120, 18091, 18091, 18091, 18067, 18067, 18067, 18038, 18038, 18038, 18014, 18014, 18014, 17985, 17985, 17985, 17961, 17961, 17961, 17932, 17932, 17932, 17908, 17908, 17908, 17879, 17879, 17855, 17855, 17855, 17826, 17826, 17826, 17802, 17802, 17802, 17772, 17772, 17772, 17749, 17749, 17749, 17719, 17719, 17719, 17696, 17696, 17696, 17666, 17666, 17666, 17642, 17642, 17642, 17613, 17613, 17613, 17589, 17589, 17560, 17560, 17560, 17536, 17536, 17536, 17506, 17506, 17506, 17483, 17483, 17483, 17453, 17453, 17453, 17429, 17429, 17429, 17400, 17400, 17400, 17376, 17376, 17376, 17346, 17346, 17346, 17323, 17323, 17323, 17293, 17293, 17269, 17269, 17269, 17240, 17240, 17240, 17216, 17216, 17216, 17186, 17186, 17186, 17162, 17162, 17162, 17133, 17133, 17133, 17109, 17109, 17109, 17079, 17079, 17079, 17055, 17055, 17055, 17026, 17026, 17026, 17002, 17002, 16972, 16972, 16972, 16948, 16948, 16948, 16925, 16925, 16925, 16895, 16895, 16895, 16871, 16871, 16871, 16841, 16841, 16841, 16817, 16817, 16817, 16788, 16788, 16788, 16764, 16764, 16764, 16734, 16734, 16734, 16710, 16710, 16680, 16680, 16680, 16657, 16657, 16657, 16627, 16627, 16627, 16603, 16603, 16603, 16573, 16573, 16573, 16549, 16549, 16549, 16519, 16519, 16519, 16495, 16495, 16495, 16465, 16465, 16465, 16442, 16442, 16442, 16412, 16412, 16388, 16388, 16388, 16358, 16358, 16358, 16334, 16334, 16334, 16304, 16304, 16304, 16280, 16280, 16280, 16250, 16250, 16250, 16226, 16226, 16226, 16196, 16196, 16196, 16172, 16172, 16172, 16142, 16142, 16142, 16118, 16118, 16118, 16088, 16088, 16064, 16064, 16064, 16034, 16034, 16034, 16010, 16010, 16010, 15980, 15980, 15980, 15956, 15956, 15956, 15926, 15926, 15926, 15902, 15902, 15902, 15872, 15872, 15872, 15848, 15848, 15848, 15818, 15818, 15818, 15794, 15794, 15794, 15764, 15764, 15740, 15740, 15740, 15716, 15716, 15716, 15686, 15686, 15686, 15662, 15662, 15662, 15632, 15632, 15632, 15608, 15608, 15608, 15577, 15577, 15577, 15553, 15553, 15553, 15523, 15523, 15523, 15499, 15499, 15499, 15469, 15469, 15469, 15445, 15445, 15415, 15415, 15415, 15391, 15391, 15391, 15360, 15360, 15360, 15336, 15336, 15336, 15306, 15306, 15306, 15282, 15282, 15282, 15252, 15252, 15252, 15227, 15227, 15227, 15197, 15197, 15197, 15173, 15173, 15173, 15143, 15143, 15143, 15119, 15119, 15088, 15088, 15088, 15064, 15064, 15064, 15034, 15034, 15034, 15010, 15010, 15010, 14979, 14979, 14979, 14955, 14955, 14955, 14925, 14925, 14925, 14900, 14900, 14900, 14870, 14870, 14870, 14846, 14846, 14846, 14816, 14816, 14816, 14791, 14791, 14791, 14761, 14761, 14737, 14737, 14737, 14706, 14706, 14706, 14682, 14682, 14682, 14652, 14652, 14652, 14627, 14627, 14627, 14597, 14597, 14597, 14572, 14572, 14572, 14542, 14542, 14542, 14518, 14518, 14518, 14493, 14493, 14493, 14463, 14463, 14463, 14439, 14439, 14439, 14408, 14408, 14384, 14384, 14384, 14353, 14353, 14353, 14329, 14329, 14329, 14298, 14298, 14298, 14274, 14274, 14274, 14243, 14243, 14243, 14219, 14219, 14219, 14188, 14188, 14188, 14164, 14164, 14164, 14133, 14133, 14133, 14109, 14109, 14109, 14078, 14078, 14078, 14054, 14054, 14023, 14023, 14023, 13999, 13999, 13999, 13968, 13968, 13968, 13944, 13944, 13944, 13913, 13913, 13913, 13889, 13889, 13889, 13858, 13858, 13858, 13834, 13834, 13834, 13803, 13803, 13803, 13778, 13778, 13778, 13748, 13748, 13748, 13723, 13723, 13723, 13693, 13693, 13693, 13668, 13668, 13637, 13637, 13637, 13613, 13613, 13613, 13582, 13582, 13582, 13557, 13557, 13557, 13527, 13527, 13527, 13502, 13502, 13502, 13471, 13471, 13471, 13447, 13447, 13447, 13416, 13416, 13416, 13391, 13391, 13391, 13361, 13361, 13361, 13336, 13336, 13336, 13305, 13305, 13305, 13280, 13280, 13256, 13256, 13256, 13225, 13225, 13225, 13200, 13200, 13200, 13169, 13169, 13169, 13145, 13145, 13145, 13114, 13114, 13114, 13089, 13089, 13089, 13058, 13058, 13058, 13034, 13034, 13034, 13003, 13003, 13003, 12978, 12978, 12978, 12947, 12947, 12947, 12922, 12922, 12922, 12891, 12891, 12891, 12867, 12867, 12836, 12836, 12836, 12811, 12811, 12811, 12780, 12780, 12780, 12755, 12755, 12755, 12724, 12724, 12724, 12699, 12699, 12699, 12668, 12668, 12668, 12643, 12643, 12643, 12612, 12612, 12612, 12588, 12588, 12588, 12557, 12557, 12557, 12532, 12532, 12532, 12501, 12501, 12501, 12476, 12476, 12476, 12445, 12445, 12445, 12420, 12420, 12389, 12389, 12389, 12364, 12364, 12364, 12333, 12333, 12333, 12308, 12308, 12308, 12277, 12277, 12277, 12252, 12252, 12252, 12221, 12221, 12221, 12196, 12196, 12196, 12164, 12164, 12164, 12139, 12139, 12139, 12108, 12108, 12108, 12083, 12083, 12083, 12058, 12058, 12058, 12027, 12027, 12027, 12002, 12002, 12002, 11971, 11971, 11946, 11946, 11946, 11915, 11915, 11915, 11890, 11890, 11890, 11858, 11858, 11858, 11833, 11833, 11833, 11802, 11802, 11802, 11777, 11777, 11777, 11746, 11746, 11746, 11721, 11721, 11721, 11689, 11689, 11689, 11664, 11664, 11664, 11633, 11633, 11633, 11608, 11608, 11608, 11576, 11576, 11576, 11551, 11551, 11551, 11520, 11520, 11520, 11495, 11495, 11463, 11463, 11463, 11438, 11438, 11438, 11407, 11407, 11407, 11382, 11382, 11382, 11350, 11350, 11350, 11325, 11325, 11325, 11293, 11293, 11293, 11268, 11268, 11268, 11237, 11237, 11237, 11212, 11212, 11212, 11180, 11180, 11180, 11155, 11155, 11155, 11123, 11123, 11123, 11098, 11098, 11098, 11067, 11067, 11067, 11041, 11041, 11041, 11010, 11010, 10984, 10984, 10984, 10953, 10953, 10953, 10928, 10928, 10928, 10896, 10896, 10896, 10871, 10871, 10871, 10839, 10839, 10839, 10814, 10814, 10814, 10788, 10788, 10788, 10757, 10757, 10757, 10731, 10731, 10731, 10700, 10700, 10700, 10674, 10674, 10674, 10643, 10643, 10643, 10617, 10617, 10617, 10586, 10586, 10586, 10560, 10560, 10560, 10528, 10528, 10528, 10503, 10503, 10503, 10471, 10471, 10446, 10446, 10446, 10414, 10414, 10414, 10389, 10389, 10389, 10357, 10357, 10357, 10331, 10331, 10331, 10300, 10300, 10300, 10274, 10274, 10274, 10242, 10242, 10242, 10217, 10217, 10217, 10185, 10185, 10185, 10159, 10159, 10159, 10128, 10128, 10128, 10102, 10102, 10102, 10070, 10070, 10070, 10045, 10045, 10045, 10013, 10013, 10013, 9987, 9987, 9987, 9955, 9955, 9955, 9930, 9930, 9930, 9898, 9898, 9898, 9872, 9872, 9840, 9840, 9840, 9814, 9814, 9814, 9782, 9782, 9782, 9757, 9757, 9757, 9725, 9725, 9725, 9699, 9699, 9699, 9667, 9667, 9667, 9641, 9641, 9641, 9609, 9609, 9609, 9584, 9584, 9584, 9552, 9552, 9552, 9526, 9526, 9526, 9500, 9500, 9500, 9468, 9468, 9468, 9442, 9442, 9442, 9410, 9410, 9410, 9385, 9385, 9385, 9352, 9352, 9352, 9327, 9327, 9327, 9294, 9294, 9294, 9269, 9269, 9269, 9236, 9236, 9236, 9211, 9211, 9178, 9178, 9178, 9153, 9153, 9153, 9120, 9120, 9120, 9095, 9095, 9095, 9062, 9062, 9062, 9036, 9036, 9036, 9004, 9004, 9004, 8978, 8978, 8978, 8946, 8946, 8946, 8920, 8920, 8920, 8888, 8888, 8888, 8862, 8862, 8862, 8830, 8830, 8830, 8804, 8804, 8804, 8771, 8771, 8771, 8745, 8745, 8745, 8713, 8713, 8713, 8687, 8687, 8687, 8655, 8655, 8655, 8629, 8629, 8629, 8596, 8596, 8596, 8570, 8570, 8570, 8538, 8538, 8538, 8512, 8512, 8512, 8479, 8479, 8453, 8453, 8453, 8421, 8421, 8421, 8395, 8395, 8395, 8362, 8362, 8362, 8336, 8336, 8336, 8303, 8303, 8303, 8277, 8277, 8277, 8245, 8245, 8245, 8219, 8219, 8219, 8193, 8193, 8193, 8160, 8160, 8160, 8134, 8134, 8134, 8101, 8101, 8101, 8075, 8075, 8075, 8042, 8042, 8042, 8016, 8016, 8016, 7984, 7984, 7984, 7957, 7957, 7957, 7925, 7925, 7925, 7899, 7899, 7899, 7866, 7866, 7866, 7840, 7840, 7840, 7807, 7807, 7807, 7781, 7781, 7781, 7748, 7748, 7748, 7722, 7722, 7722, 7689, 7689, 7689, 7663, 7663, 7663, 7630, 7630, 7630, 7603, 7603, 7571, 7571, 7571, 7544, 7544, 7544, 7511, 7511, 7511, 7485, 7485, 7485, 7452, 7452, 7452, 7426, 7426, 7426, 7393, 7393, 7393, 7367, 7367, 7367, 7334, 7334, 7334, 7307, 7307, 7307, 7274, 7274, 7274, 7248, 7248, 7248, 7215, 7215, 7215, 7188, 7188, 7188, 7155, 7155, 7155, 7129, 7129, 7129, 7096, 7096, 7096, 7070, 7070, 7070, 7036, 7036, 7036, 7010, 7010, 7010, 6977, 6977, 6977, 6950, 6950, 6950, 6924, 6924, 6924, 6891, 6891, 6891, 6864, 6864, 6864, 6831, 6831, 6831, 6805, 6805, 6805, 6771, 6771, 6771, 6745, 6745, 6745, 6712, 6712, 6712, 6685, 6685, 6685, 6652, 6652, 6652, 6625, 6625, 6625, 6592, 6592, 6592, 6565, 6565, 6565, 6532, 6532, 6532, 6506, 6506, 6506, 6472, 6472, 6446, 6446, 6446, 6412, 6412, 6412, 6386, 6386, 6386, 6352, 6352, 6352, 6326, 6326, 6326, 6292, 6292, 6292, 6265, 6265, 6265, 6232, 6232, 6232, 6205, 6205, 6205, 6172, 6172, 6172, 6145, 6145, 6145, 6112, 6112, 6112, 6085, 6085, 6085, 6051, 6051, 6051, 6025, 6025, 6025, 5991, 5991, 5991, 5964, 5964, 5964, 5931, 5931, 5931, 5904, 5904, 5904, 5870, 5870, 5870, 5844, 5844, 5844, 5810, 5810, 5810, 5783, 5783, 5783, 5750, 5750, 5750, 5723, 5723, 5723, 5689, 5689, 5689, 5662, 5662, 5662, 5628, 5628, 5628, 5601, 5601, 5601, 5575, 5575, 5575, 5541, 5541, 5541, 5514, 5514, 5514, 5480, 5480, 5480, 5453, 5453, 5453, 5419, 5419, 5419, 5392, 5392, 5392, 5359, 5359, 5359, 5332, 5332, 5332, 5298, 5298, 5298, 5271, 5271, 5271, 5237, 5237, 5237, 5210, 5210, 5210, 5176, 5176, 5176, 5149, 5149, 5149, 5115, 5115, 5115, 5088, 5088, 5088, 5054, 5054, 5054, 5027, 5027, 5027, 4993, 4993, 4993, 4966, 4966, 4966, 4932, 4932, 4932, 4905, 4905, 4905, 4871, 4871, 4871, 4844, 4844, 4844, 4810, 4810, 4810, 4782, 4782, 4782, 4748, 4748, 4748, 4721, 4721, 4721, 4687, 4687, 4687, 4660, 4660, 4660, 4626, 4626, 4626, 4598, 4598, 4598, 4564, 4564, 4564, 4537, 4537, 4537, 4503, 4503, 4503, 4475, 4475, 4475, 4441, 4441, 4441, 4414, 4414, 4414, 4380, 4380, 4380, 4352, 4352, 4352, 4318, 4318, 4318, 4291, 4291, 4291, 4257, 4257, 4257, 4229, 4229, 4229, 4202, 4202, 4202, 4167, 4167, 4167, 4140, 4140, 4140, 4106, 4106, 4106, 4078, 4078, 4078, 4044, 4044, 4016, 4016, 4016, 3982, 3982, 3982, 3954, 3954, 3954, 3920, 3920, 3920, 3893, 3893, 3893, 3858, 3858, 3858, 3831, 3831, 3831, 3796, 3796, 3796, 3769, 3769, 3769, 3734, 3734, 3734, 3706, 3706, 3706, 3672, 3672, 3672, 3644, 3644, 3644, 3610, 3610, 3610, 3582, 3582, 3582, 3548, 3548, 3548, 3520, 3520, 3520, 3485, 3485, 3485, 3458, 3458, 3458, 3423, 3423, 3423, 3395, 3395, 3395, 3361, 3361, 3361, 3333, 3333, 3333, 3298, 3298, 3298, 3298, 3270, 3270, 3270, 3236, 3236, 3236, 3208, 3208, 3208, 3173, 3173, 3173, 3145, 3145, 3145, 3111, 3111, 3111, 3083, 3083, 3083, 3048, 3048, 3048, 3020, 3020, 3020, 2985, 2985, 2985, 2957, 2957, 2957, 2923, 2923, 2923, 2895, 2895, 2895, 2860, 2860, 2860, 2832, 2832, 2832, 2804, 2804, 2804, 2769, 2769, 2769, 2741, 2741, 2741, 2706, 2706, 2706, 2678, 2678, 2678, 2643, 2643, 2643, 2615, 2615, 2615, 2580, 2580, 2580, 2552, 2552, 2552, 2517, 2517, 2517, 2489, 2489, 2489, 2454, 2454, 2454, 2426, 2426, 2426, 2391, 2391, 2391, 2363, 2363, 2363, 2328, 2328, 2328, 2299, 2299, 2299, 2264, 2264, 2264, 2236, 2236, 2236, 2201, 2201, 2201, 2173, 2173, 2173, 2138, 2138, 2138, 2109, 2109, 2109, 2074, 2074, 2074, 2046, 2046, 2046, 2011, 2011, 2011, 1982, 1982, 1982, 1947, 1947, 1947, 1919, 1919, 1919, 1883, 1883, 1883, 1855, 1855, 1855, 1820, 1820, 1820, 1792, 1792, 1792, 1756, 1756, 1756, 1728, 1728, 1728, 1692, 1692, 1692, 1664, 1664, 1664, 1629, 1629, 1629, 1600, 1600, 1600, 1565, 1565, 1565, 1536, 1536, 1536, 1501, 1501, 1501, 1472, 1472, 1472, 1437, 1437, 1437, 1408, 1408, 1408, 1380, 1380, 1380, 1344, 1344, 1344, 1316, 1316, 1316, 1280, 1280, 1280, 1252, 1252, 1252, 1216, 1216, 1216, 1187, 1187, 1187, 1152, 1152, 1152, 1123, 1123, 1123, 1087, 1087, 1087, 1059, 1059, 1059, 1023, 1023, 1023, 994, 994, 994, 959, 959, 959, 930, 930, 930, 894, 894, 894, 894, 865, 865, 865, 830, 830, 830, 801, 801, 801, 765, 765, 765, 736, 736, 736, 700, 700, 700, 672, 672, 672, 636, 636, 636, 607, 607, 607, 571, 571, 571, 542, 542, 542, 506, 506, 506, 477, 477, 477, 441, 441, 441, 412, 412, 412, 376, 376, 376, 347, 347, 347, 311, 311, 311, 282, 282, 282, 246, 246, 246, 217, 217, 217, 181, 181, 181, 152, 152, 152, 116, 116, 116, 87, 87, 87, 51, 51, 51, 22, 22, 22, 71993, 71993, 71993, 71956, 71956, 71956, 71927, 71927, 71927, 71891, 71891, 71891, 71862, 71862, 71862, 71826, 71826, 71826, 71797, 71797, 71797, 71761, 71761, 71761, 71732, 71732, 71732, 71732, 71696, 71696, 71696, 71667, 71667, 71667, 71631, 71631, 71631, 71602, 71602, 71602, 71566, 71566, 71566, 71537, 71537, 71537, 71501, 71501, 71501, 71472, 71472, 71472, 71436, 71436, 71436, 71408, 71408, 71408, 71372, 71372, 71372, 71343, 71343, 71343, 71307, 71307, 71307, 71278, 71278, 71278, 71242, 71242, 71242, 71213, 71213, 71213, 71178, 71178, 71178, 71149, 71149, 71149, 71113, 71113, 71113, 71084, 71084, 71084, 71049, 71049, 71049, 71020, 71020, 71020, 70984, 70984, 70984, 70956, 70956, 70956, 70920, 70920, 70920, 70891, 70891, 70891, 70856, 70856, 70856, 70856, 70827, 70827, 70827, 70791, 70791, 70791, 70763, 70763, 70763, 70727, 70727, 70727, 70699, 70699, 70699, 70663, 70663, 70663, 70634, 70634, 70634, 70599, 70599, 70599, 70570, 70570, 70570, 70542, 70542, 70542, 70506, 70506, 70506, 70478, 70478, 70478, 70442, 70442, 70442, 70414, 70414, 70414, 70379, 70379, 70379, 70350, 70350, 70350, 70315, 70315, 70315, 70286, 70286, 70286, 70251, 70251, 70251, 70223, 70223, 70223, 70187, 70187, 70187, 70159, 70159, 70159, 70159, 70124, 70124, 70124, 70095, 70095, 70095, 70060, 70060, 70060, 70032, 70032, 70032, 69996, 69996, 69996, 69968, 69968, 69968, 69933, 69933, 69933, 69905, 69905, 69905, 69869, 69869, 69869, 69841, 69841, 69841, 69806, 69806, 69806, 69778, 69778, 69778, 69743, 69743, 69743, 69715, 69715, 69715, 69679, 69679, 69679, 69651, 69651, 69651, 69616, 69616, 69616, 69588, 69588, 69588, 69553, 69553, 69553, 69525, 69525, 69525, 69525, 69490, 69490, 69490, 69462, 69462, 69462, 69427, 69427, 69427, 69399, 69399, 69399, 69364, 69364, 69364, 69336, 69336, 69336, 69301, 69301, 69301, 69273, 69273, 69273, 69238, 69238, 69238, 69210, 69210, 69210, 69175, 69175, 69175, 69147, 69147, 69147, 69119, 69119, 69119, 69084, 69084, 69084, 69056, 69056, 69056, 69022, 69022, 69022, 68994, 68994, 68994, 68959, 68959, 68959, 68959, 68931, 68931, 68931, 68896, 68896, 68896, 68868, 68868, 68868, 68834, 68834, 68834, 68806, 68806, 68806, 68771, 68771, 68771, 68743, 68743, 68743, 68709, 68709, 68709, 68681, 68681, 68681, 68646, 68646, 68646, 68619, 68619, 68619, 68584, 68584, 68584, 68556, 68556, 68556, 68522, 68522, 68522, 68494, 68494, 68494, 68459, 68459, 68459, 68459, 68432, 68432, 68432, 68397, 68397, 68397, 68369, 68369, 68369, 68335, 68335, 68335, 68307, 68307, 68307, 68273, 68273, 68273, 68245, 68245, 68245, 68211, 68211, 68211, 68183, 68183, 68183, 68149, 68149, 68149, 68121, 68121, 68121, 68087, 68087, 68087, 68059, 68059, 68059, 68025, 68025, 68025, 67997, 67997, 67997, 67997, 67963, 67963, 67963, 67936, 67936, 67936, 67901, 67901, 67901, 67874, 67874, 67874, 67839, 67839, 67839, 67812, 67812, 67812, 67778, 67778, 67778, 67750, 67750, 67750, 67723, 67723, 67723, 67689, 67689, 67689, 67661, 67661, 67661, 67627, 67627, 67627, 67600, 67600, 67600, 67566, 67566, 67566, 67566, 67538, 67538, 67538, 67504, 67504, 67504, 67477, 67477, 67477, 67443, 67443, 67443, 67415, 67415, 67415, 67381, 67381, 67381, 67354, 67354, 67354, 67320, 67320, 67320, 67293, 67293, 67293, 67259, 67259, 67259, 67231, 67231, 67231, 67197, 67197, 67197, 67170, 67170, 67170, 67170, 67136, 67136, 67136, 67109, 67109, 67109, 67075, 67075, 67075, 67048, 67048, 67048, 67014, 67014, 67014, 66987, 66987, 66987, 66953, 66953, 66953, 66926, 66926, 66926, 66892, 66892, 66892, 66865, 66865, 66865, 66831, 66831, 66831, 66804, 66804, 66804, 66804, 66770, 66770, 66770, 66743, 66743, 66743, 66709, 66709, 66709, 66682, 66682, 66682, 66648, 66648, 66648, 66621, 66621, 66621, 66587, 66587, 66587, 66560, 66560, 66560, 66527, 66527, 66527, 66500, 66500, 66500, 66466, 66466, 66466, 66439, 66439, 66439, 66439, 66412, 66412, 66412, 66378, 66378, 66378, 66351, 66351, 66351, 66318, 66318, 66318, 66291, 66291, 66291, 66257, 66257, 66257, 66230, 66230, 66230, 66197, 66197, 66197, 66170, 66170, 66170, 66136, 66136, 66136, 66109, 66109, 66109, 66076, 66076, 66076, 66076, 66049, 66049, 66049, 66016, 66016, 66016, 65989, 65989, 65989, 65955, 65955, 65955, 65928, 65928, 65928, 65895, 65895, 65895, 65868, 65868, 65868, 65835, 65835, 65835, 65808, 65808, 65808, 65775, 65775, 65775, 65748, 65748, 65748, 65748, 65715, 65715, 65715, 65688, 65688, 65688, 65654, 65654, 65654, 65628, 65628, 65628, 65594, 65594, 65594, 65568, 65568, 65568, 65534, 65534, 65534, 65508, 65508, 65508, 65475, 65475, 65475, 65448, 65448, 65448, 65448, 65415, 65415, 65415, 65388, 65388, 65388, 65355, 65355, 65355, 65328, 65328, 65328, 65295, 65295, 65295, 65268, 65268, 65268, 65235, 65235, 65235, 65209, 65209, 65209, 65175, 65175, 65175, 65149, 65149, 65149, 65149, 65116, 65116, 65116, 65089, 65089, 65089, 65063, 65063, 65063, 65030, 65030, 65030, 65003, 65003, 65003, 64970, 64970, 64970, 64944, 64944, 64944, 64911, 64911, 64911, 64884, 64884, 64884, 64851, 64851, 64851, 64851, 64825, 64825, 64825, 64792, 64792, 64792, 64765, 64765, 64765, 64732, 64732, 64732, 64706, 64706, 64706, 64673, 64673, 64673, 64647, 64647, 64647, 64614, 64614, 64614, 64587, 64587, 64587, 64587, 64554, 64554, 64554, 64528, 64528, 64528, 64495, 64495, 64495, 64469, 64469, 64469, 64436, 64436, 64436, 64410, 64410, 64410, 64377, 64377, 64377, 64351, 64351, 64351, 64318, 64318, 64318, 64318, 64292, 64292, 64292, 64259, 64259, 64259, 64232, 64232, 64232, 64200, 64200, 64200, 64173, 64173, 64173, 64141, 64141, 64141, 64115, 64115, 64115, 64082, 64082, 64082, 64056, 64056, 64056, 64056, 64023, 64023, 64023, 63997, 63997, 63997, 63964, 63964, 63964, 63938, 63938, 63938, 63905, 63905, 63905, 63879, 63879, 63879, 63847, 63847, 63847, 63820, 63820, 63820, 63788, 63788, 63788, 63788, 63762, 63762, 63762, 63736, 63736, 63736, 63703, 63703, 63703, 63677, 63677, 63677, 63644, 63644, 63644, 63618, 63618, 63618, 63586, 63586, 63586, 63560, 63560, 63560, 63560, 63527, 63527, 63527, 63501, 63501, 63501, 63469, 63469, 63469, 63443, 63443, 63443, 63410, 63410, 63410, 63384, 63384, 63384, 63352, 63352, 63352, 63326, 63326, 63326, 63326, 63294, 63294, 63294, 63268, 63268, 63268, 63235, 63235, 63235, 63209, 63209, 63209, 63177, 63177, 63177, 63151, 63151, 63151, 63119, 63119, 63119, 63093, 63093, 63093, 63093, 63060, 63060, 63060, 63035, 63035, 63035, 63002, 63002, 63002, 62976, 62976, 62976, 62944, 62944, 62944, 62918, 62918, 62918, 62886, 62886, 62886, 62860, 62860, 62860, 62860, 62828, 62828, 62828, 62802, 62802, 62802, 62770, 62770, 62770, 62744, 62744, 62744, 62712, 62712, 62712, 62686, 62686, 62686, 62654, 62654, 62654, 62628, 62628, 62628, 62628, 62596, 62596, 62596, 62570, 62570, 62570, 62538, 62538, 62538, 62513, 62513, 62513, 62480, 62480, 62480, 62455, 62455, 62455, 62429, 62429, 62429, 62429, 62397, 62397, 62397, 62371, 62371, 62371, 62339, 62339, 62339, 62314, 62314, 62314, 62282, 62282, 62282, 62256, 62256, 62256, 62224, 62224, 62224, 62198, 62198, 62198, 62198, 62166, 62166, 62166, 62141, 62141, 62141, 62109, 62109, 62109, 62083, 62083, 62083, 62051, 62051, 62051, 62026, 62026, 62026, 61994, 61994, 61994, 61994, 61968, 61968, 61968, 61936, 61936, 61936, 61911, 61911, 61911, 61879, 61879, 61879, 61853, 61853, 61853, 61821, 61821, 61821, 61796, 61796, 61796, 61796, 61764, 61764, 61764, 61739, 61739, 61739, 61707, 61707, 61707, 61681, 61681, 61681, 61649, 61649, 61649, 61624, 61624, 61624, 61592, 61592, 61592, 61592, 61567, 61567, 61567, 61535, 61535, 61535, 61510, 61510, 61510, 61478, 61478, 61478, 61452, 61452, 61452, 61421, 61421, 61421, 61421, 61395, 61395, 61395, 61364, 61364, 61364, 61338, 61338, 61338, 61307, 61307, 61307, 61281, 61281, 61281, 61250, 61250, 61250, 61224, 61224, 61224, 61224, 61193, 61193, 61193, 61167, 61167, 61167, 61142, 61142, 61142, 61110, 61110, 61110, 61085, 61085, 61085, 61053, 61053, 61053, 61028, 61028, 61028, 61028, 60997, 60997, 60997, 60971, 60971, 60971, 60940, 60940, 60940, 60915, 60915, 60915, 60883, 60883, 60883, 60858, 60858, 60858, 60858, 60826, 60826, 60826, 60801, 60801, 60801, 60769, 60769, 60769, 60744, 60744, 60744, 60713, 60713, 60713, 60688, 60688, 60688, 60688, 60656, 60656, 60656, 60631, 60631, 60631, 60600, 60600, 60600, 60574, 60574, 60574, 60543, 60543, 60543, 60518, 60518, 60518, 60486, 60486, 60486, 60486, 60461, 60461, 60461, 60430, 60430, 60430, 60405, 60405, 60405, 60373, 60373, 60373, 60348, 60348, 60348, 60317, 60317, 60317, 60317, 60292, 60292, 60292, 60261, 60261, 60261, 60236, 60236, 60236, 60204, 60204, 60204, 60179, 60179, 60179, 60148, 60148, 60148, 60148, 60123, 60123, 60123, 60092, 60092, 60092, 60067, 60067, 60067, 60035, 60035, 60035, 60010, 60010, 60010, 59979, 59979, 59979, 59979, 59954, 59954, 59954, 59929, 59929, 59929, 59898, 59898, 59898, 59873, 59873, 59873, 59842, 59842, 59842, 59842, 59817, 59817, 59817, 59786, 59786, 59786, 59761, 59761, 59761, 59730, 59730, 59730, 59705, 59705, 59705, 59674, 59674, 59674, 59674, 59649, 59649, 59649, 59618, 59618, 59618, 59593, 59593, 59593, 59562, 59562, 59562, 59537, 59537, 59537, 59506, 59506, 59506, 59506, 59481, 59481, 59481, 59450, 59450, 59450, 59425, 59425, 59425, 59394, 59394, 59394, 59369, 59369, 59369, 59369, 59338, 59338, 59338, 59313, 59313, 59313, 59282, 59282, 59282, 59257, 59257, 59257, 59226, 59226, 59226, 59202, 59202, 59202, 59202, 59171, 59171, 59171, 59146, 59146, 59146, 59115, 59115, 59115, 59090, 59090, 59090, 59059, 59059, 59059, 59059, 59034, 59034, 59034, 59004, 59004, 59004, 58979, 58979, 58979, 58948, 58948, 58948, 58923, 58923, 58923, 58892, 58892, 58892, 58892, 58868, 58868, 58868, 58837, 58837, 58837, 58812, 58812, 58812, 58781, 58781, 58781, 58757, 58757, 58757, 58757, 58726, 58726, 58726, 58701, 58701, 58701, 58676, 58676, 58676, 58646, 58646, 58646, 58621, 58621, 58621, 58621, 58590, 58590, 58590, 58566, 58566, 58566, 58535, 58535, 58535, 58510, 58510, 58510, 58479, 58479, 58479, 58455, 58455, 58455, 58455, 58424, 58424, 58424, 58400, 58400, 58400, 58369, 58369, 58369, 58344, 58344, 58344, 58314, 58314, 58314, 58314, 58289, 58289, 58289, 58258, 58258, 58258, 58234, 58234, 58234, 58203, 58203, 58203, 58179, 58179, 58179, 58179, 58148, 58148, 58148, 58124, 58124, 58124, 58093, 58093, 58093, 58068, 58068, 58068, 58038, 58038, 58038, 58038, 58013, 58013, 58013, 57983, 57983, 57983, 57958, 57958, 57958, 57928, 57928, 57928, 57903, 57903, 57903, 57903, 57873, 57873, 57873, 57848, 57848, 57848, 57818, 57818, 57818, 57793, 57793, 57793, 57763, 57763, 57763, 57763, 57738, 57738, 57738, 57708, 57708, 57708, 57683, 57683, 57683, 57653, 57653, 57653, 57629, 57629, 57629, 57629, 57598, 57598, 57598, 57574, 57574, 57574, 57543, 57543, 57543, 57519, 57519, 57519, 57519, 57488, 57488, 57488, 57464, 57464, 57464, 57440, 57440, 57440, 57409, 57409, 57409, 57385, 57385, 57385, 57385, 57355, 57355, 57355, 57330, 57330, 57330, 57300, 57300, 57300, 57276, 57276, 57276, 57245, 57245, 57245, 57245, 57221, 57221, 57221, 57191, 57191, 57191, 57166, 57166, 57166, 57136, 57136, 57136, 57136, 57112, 57112, 57112, 57081, 57081, 57081, 57057, 57057, 57057, 57027, 57027, 57027, 57003, 57003, 57003, 57003, 56972, 56972, 56972, 56948, 56948, 56948, 56918, 56918, 56918, 56894, 56894, 56894, 56863, 56863, 56863, 56863, 56839, 56839, 56839, 56809, 56809, 56809, 56785, 56785, 56785, 56754, 56754, 56754, 56754, 56730, 56730, 56730, 56700, 56700, 56700, 56676, 56676, 56676, 56646, 56646, 56646, 56622, 56622, 56622, 56622, 56591, 56591, 56591, 56567, 56567, 56567, 56537, 56537, 56537, 56513, 56513, 56513, 56513, 56483, 56483, 56483, 56459, 56459, 56459, 56429, 56429, 56429, 56404, 56404, 56404, 56404, 56374, 56374, 56374, 56350, 56350, 56350, 56320, 56320, 56320, 56296, 56296, 56296, 56266, 56266, 56266, 56266, 56242, 56242, 56242, 56218, 56218, 56218, 56188, 56188, 56188, 56164, 56164, 56164, 56164, 56134, 56134, 56134, 56110, 56110, 56110, 56080, 56080, 56080, 56056, 56056, 56056, 56056, 56026, 56026, 56026, 56002, 56002, 56002, 55972, 55972, 55972, 55948, 55948, 55948, 55918, 55918, 55918, 55918, 55894, 55894, 55894, 55864, 55864, 55864, 55840, 55840, 55840, 55810, 55810, 55810, 55810, 55786, 55786, 55786, 55756, 55756, 55756, 55732, 55732, 55732, 55702, 55702, 55702, 55702, 55678, 55678, 55678, 55648, 55648, 55648, 55624, 55624, 55624, 55594, 55594, 55594, 55594, 55570, 55570, 55570, 55541, 55541, 55541, 55517, 55517, 55517, 55487, 55487, 55487, 55487, 55463, 55463, 55463, 55433, 55433, 55433, 55409, 55409, 55409, 55379, 55379, 55379, 55379, 55355, 55355, 55355, 55326, 55326, 55326, 55302, 55302, 55302, 55272, 55272, 55272, 55272, 55248, 55248, 55248, 55218, 55218, 55218, 55194, 55194, 55194, 55165, 55165, 55165, 55165, 55141, 55141, 55141, 55111, 55111, 55111, 55087, 55087, 55087, 55063, 55063, 55063, 55063, 55034, 55034, 55034, 55010, 55010, 55010, 54980, 54980, 54980, 54956, 54956, 54956, 54956, 54927, 54927, 54927, 54903, 54903, 54903, 54873, 54873, 54873, 54849, 54849, 54849, 54849, 54820, 54820, 54820, 54796, 54796, 54796, 54766, 54766, 54766, 54743, 54743, 54743, 54743, 54713, 54713, 54713, 54689, 54689, 54689, 54660, 54660, 54660, 54636, 54636, 54636, 54636, 54606, 54606, 54606, 54583, 54583, 54583, 54553, 54553, 54553, 54529, 54529, 54529, 54529, 54500, 54500, 54500, 54476, 54476, 54476, 54446, 54446, 54446, 54446, 54423, 54423, 54423, 54393, 54393, 54393, 54369, 54369, 54369, 54340, 54340, 54340, 54340, 54316, 54316, 54316, 54287, 54287, 54287, 54263, 54263, 54263, 54234, 54234, 54234, 54234, 54210, 54210, 54210, 54180, 54180, 54180, 54157, 54157, 54157, 54127, 54127, 54127, 54127, 54104, 54104, 54104, 54074, 54074, 54074, 54051, 54051, 54051, 54051, 54021, 54021, 54021, 53998, 53998, 53998, 53968, 53968, 53968, 53944, 53944, 53944, 53944, 53915, 53915, 53915, 53891, 53891, 53891, 53868, 53868, 53868, 53838, 53838, 53838, 53838, 53815, 53815, 53815, 53785, 53785, 53785, 53762, 53762, 53762, 53762, 53733, 53733, 53733, 53709, 53709, 53709, 53680, 53680, 53680, 53656, 53656, 53656, 53656, 53627, 53627, 53627, 53603, 53603, 53603, 53574, 53574, 53574, 53574, 53550, 53550, 53550, 53521, 53521, 53521, 53498, 53498, 53498, 53468, 53468, 53468, 53468, 53445, 53445, 53445, 53415, 53415, 53415, 53392, 53392, 53392, 53392, 53363, 53363, 53363, 53339, 53339, 53339, 53310, 53310, 53310, 53286, 53286, 53286, 53286, 53257, 53257, 53257, 53234, 53234, 53234, 53204, 53204, 53204, 53204, 53181, 53181, 53181, 53152, 53152, 53152, 53128, 53128, 53128, 53099, 53099, 53099, 53099, 53076, 53076, 53076, 53046, 53046, 53046, 53023, 53023, 53023, 53023, 52994, 52994, 52994, 52970, 52970, 52970, 52941, 52941, 52941, 52918, 52918, 52918, 52918, 52889, 52889, 52889, 52865, 52865, 52865, 52836, 52836, 52836, 52836, 52813, 52813, 52813, 52783, 52783, 52783, 52760, 52760, 52760, 52760, 52731, 52731, 52731, 52708, 52708, 52708, 52684, 52684, 52684, 52655, 52655, 52655, 52655, 52632, 52632, 52632, 52603, 52603, 52603, 52579, 52579, 52579, 52579, 52550, 52550, 52550, 52527, 52527, 52527, 52498, 52498, 52498, 52498, 52475, 52475, 52475, 52445, 52445, 52445, 52422, 52422, 52422, 52393, 52393, 52393, 52393, 52370, 52370, 52370, 52341, 52341, 52341, 52318, 52318, 52318, 52318, 52288, 52288, 52288, 52265, 52265, 52265, 52236, 52236, 52236, 52236, 52213, 52213, 52213, 52184, 52184, 52184, 52161, 52161, 52161, 52161, 52132, 52132, 52132, 52108, 52108, 52108, 52079, 52079, 52079, 52079, 52056, 52056, 52056, 52027, 52027, 52027, 52004, 52004, 52004, 51975, 51975, 51975, 51975, 51952, 51952, 51952, 51923, 51923, 51923, 51900, 51900, 51900, 51900, 51871, 51871, 51871, 51847, 51847, 51847, 51818, 51818, 51818, 51818, 51795, 51795, 51795, 51766, 51766, 51766, 51743, 51743, 51743, 51743, 51714, 51714, 51714, 51691, 51691, 51691, 51662, 51662, 51662, 51662, 51639, 51639, 51639, 51610, 51610, 51610, 51587, 51587, 51587, 51587, 51558, 51558, 51558, 51535, 51535, 51535, 51512, 51512, 51512, 51512, 51483, 51483, 51483, 51460, 51460, 51460, 51431, 51431, 51431, 51431, 51408, 51408, 51408, 51379, 51379, 51379, 51356, 51356, 51356, 51356, 51327, 51327, 51327, 51304, 51304, 51304, 51275, 51275, 51275, 51252, 51252, 51252, 51252, 51223, 51223, 51223, 51200, 51200, 51200, 51171, 51171, 51171, 51171, 51148, 51148, 51148, 51120, 51120, 51120, 51096, 51096, 51096, 51096, 51068, 51068, 51068, 51045, 51045, 51045, 51016, 51016, 51016, 51016, 50993, 50993, 50993, 50964, 50964, 50964, 50964, 50941, 50941, 50941, 50912, 50912, 50912, 50889, 50889, 50889, 50889, 50861, 50861, 50861, 50838, 50838, 50838, 50809, 50809, 50809, 50809, 50786, 50786, 50786, 50757, 50757, 50757, 50734, 50734, 50734, 50734, 50705, 50705, 50705, 50682, 50682, 50682, 50654, 50654, 50654, 50654, 50631, 50631, 50631, 50602, 50602, 50602, 50579, 50579, 50579, 50579, 50550, 50550, 50550, 50527, 50527, 50527, 50499, 50499, 50499, 50499, 50476, 50476, 50476, 50447, 50447, 50447, 50424, 50424, 50424, 50424, 50396, 50396, 50396, 50373, 50373, 50373, 50350, 50350, 50350, 50350, 50321, 50321, 50321, 50298, 50298, 50298, 50269, 50269, 50269, 50269, 50247, 50247, 50247, 50218, 50218, 50218, 50218, 50195, 50195, 50195, 50166, 50166, 50166, 50144, 50144, 50144, 50144, 50115, 50115, 50115, 50092, 50092, 50092, 50063, 50063, 50063, 50063, 50041, 50041, 50041, 50012, 50012, 50012, 49989, 49989, 49989, 49989, 49961, 49961, 49961, 49938, 49938, 49938, 49938, 49909, 49909, 49909, 49886, 49886, 49886, 49858, 49858, 49858, 49858, 49835, 49835, 49835, 49806, 49806, 49806, 49784, 49784, 49784, 49784, 49755, 49755, 49755, 49732, 49732, 49732, 49704, 49704, 49704, 49704, 49681, 49681, 49681, 49652, 49652, 49652, 49652, 49630, 49630, 49630, 49601, 49601, 49601, 49578, 49578, 49578, 49578, 49550, 49550, 49550, 49527, 49527, 49527, 49498, 49498, 49498, 49498, 49476, 49476, 49476, 49447, 49447, 49447, 49424, 49424, 49424, 49424, 49396, 49396, 49396, 49373, 49373, 49373, 49373, 49345, 49345, 49345, 49322, 49322, 49322, 49294, 49294, 49294, 49294, 49271, 49271, 49271, 49248, 49248, 49248, 49248, 49220, 49220, 49220, 49197, 49197, 49197, 49168, 49168, 49168, 49168, 49146, 49146, 49146, 49117, 49117, 49117, 49095, 49095, 49095, 49095, 49066, 49066, 49066, 49043, 49043, 49043, 49043, 49015, 49015, 49015, 48992, 48992, 48992, 48964, 48964, 48964, 48964, 48941, 48941, 48941, 48913, 48913, 48913, 48890, 48890, 48890, 48890, 48862, 48862, 48862, 48839, 48839, 48839, 48839, 48811, 48811, 48811, 48788, 48788, 48788, 48760, 48760, 48760, 48760, 48737, 48737, 48737, 48709, 48709, 48709, 48709, 48686, 48686, 48686, 48658, 48658, 48658, 48635, 48635, 48635, 48635, 48607, 48607, 48607, 48584, 48584, 48584, 48584, 48556, 48556, 48556, 48533, 48533, 48533, 48505, 48505, 48505, 48505, 48482, 48482, 48482, 48454, 48454, 48454, 48454, 48431, 48431, 48431, 48403, 48403, 48403, 48380, 48380, 48380, 48380, 48352, 48352, 48352, 48329, 48329, 48329, 48329, 48301, 48301, 48301, 48279, 48279, 48279, 48250, 48250, 48250, 48250, 48228, 48228, 48228, 48199, 48199, 48199, 48199, 48177, 48177, 48177, 48149, 48149, 48149, 48126, 48126, 48126, 48126, 48103, 48103, 48103, 48075, 48075, 48075, 48075, 48053, 48053, 48053, 48024, 48024, 48024, 48002, 48002, 48002, 48002, 47974, 47974, 47974, 47951, 47951, 47951, 47951, 47923, 47923, 47923, 47900, 47900, 47900, 47872, 47872, 47872, 47872, 47850, 47850, 47850, 47821, 47821, 47821, 47821, 47799, 47799, 47799, 47771, 47771, 47771, 47771, 47748, 47748, 47748, 47720, 47720, 47720, 47697, 47697, 47697, 47697, 47669, 47669, 47669, 47647, 47647, 47647, 47647, 47619, 47619, 47619, 47596, 47596, 47596, 47568, 47568, 47568, 47568, 47545, 47545, 47545, 47517, 47517, 47517, 47517, 47495, 47495, 47495, 47467, 47467, 47467, 47467, 47444, 47444, 47444, 47416, 47416, 47416, 47393, 47393, 47393, 47393, 47365, 47365, 47365, 47343, 47343, 47343, 47343, 47315, 47315, 47315, 47292, 47292, 47292, 47292, 47264, 47264, 47264, 47242, 47242, 47242, 47214, 47214, 47214, 47214, 47191, 47191, 47191, 47163, 47163, 47163, 47163, 47141, 47141, 47141, 47113, 47113, 47113, 47113, 47090, 47090, 47090, 47062, 47062, 47062, 47040, 47040, 47040, 47040, 47011, 47011, 47011, 46989, 46989, 46989, 46989, 46967, 46967, 46967, 46939, 46939, 46939, 46939, 46916, 46916, 46916, 46888, 46888, 46888, 46888, 46866, 46866, 46866, 46838, 46838, 46838, 46815, 46815, 46815, 46815, 46787, 46787, 46787, 46765, 46765, 46765, 46765, 46737, 46737, 46737, 46714, 46714, 46714, 46714, 46686, 46686, 46686, 46664, 46664, 46664, 46664, 46636, 46636, 46636, 46614, 46614, 46614, 46586, 46586, 46586, 46586, 46563, 46563, 46563, 46535, 46535, 46535, 46535, 46513, 46513, 46513, 46485, 46485, 46485, 46485, 46462, 46462, 46462, 46434, 46434, 46434, 46434, 46412, 46412, 46412, 46384, 46384, 46384, 46362, 46362, 46362, 46362, 46334, 46334, 46334, 46311, 46311, 46311, 46311, 46283, 46283, 46283, 46261, 46261, 46261, 46261, 46233, 46233, 46233, 46211, 46211, 46211, 46211, 46183, 46183, 46183, 46161, 46161, 46161, 46161, 46133, 46133, 46133, 46110, 46110, 46110, 46110, 46082, 46082, 46082, 46060, 46060, 46060, 46032, 46032, 46032, 46032, 46010, 46010, 46010, 45982, 45982, 45982, 45982, 45960, 45960, 45960, 45932, 45932, 45932, 45932, 45909, 45909, 45909, 45881, 45881, 45881, 45881, 45859, 45859, 45859, 45837, 45837, 45837, 45837, 45809, 45809, 45809, 45787, 45787, 45787, 45787, 45759, 45759, 45759, 45736, 45736, 45736, 45736, 45709, 45709, 45709, 45686, 45686, 45686, 45658, 45658, 45658, 45658, 45636, 45636, 45636, 45608, 45608, 45608, 45608, 45586, 45586, 45586, 45558, 45558, 45558, 45558, 45536, 45536, 45536, 45508, 45508, 45508, 45508, 45486, 45486, 45486, 45458, 45458, 45458, 45458, 45436, 45436, 45436, 45408, 45408, 45408, 45408, 45386, 45386, 45386, 45358, 45358, 45358, 45358, 45336, 45336, 45336, 45308, 45308, 45308, 45308, 45285, 45285, 45285, 45258, 45258, 45258, 45258, 45235, 45235, 45235, 45208, 45208, 45208, 45208, 45185, 45185, 45185, 45158, 45158, 45158, 45158, 45135, 45135, 45135, 45108, 45108, 45108, 45108, 45085, 45085, 45085, 45058, 45058, 45058, 45058, 45035, 45035, 45035, 45008, 45008, 45008, 45008, 44985, 44985, 44985, 44958, 44958, 44958, 44958, 44935, 44935, 44935, 44908, 44908, 44908, 44908, 44885, 44885, 44885, 44858, 44858, 44858, 44858, 44835, 44835, 44835, 44808, 44808, 44808, 44808, 44785, 44785, 44785, 44763, 44763, 44763, 44763, 44736, 44736, 44736, 44713, 44713, 44713, 44713, 44686, 44686, 44686, 44663, 44663, 44663, 44663, 44636, 44636, 44636, 44613, 44613, 44613, 44613, 44586, 44586, 44586, 44564, 44564, 44564, 44564, 44536, 44536, 44536, 44514, 44514, 44514, 44514, 44486, 44486, 44486, 44464, 44464, 44464, 44464, 44436, 44436, 44436, 44414, 44414, 44414, 44414, 44386, 44386, 44386, 44364, 44364, 44364, 44364, 44336, 44336, 44336, 44314, 44314, 44314, 44314, 44287, 44287, 44287, 44264, 44264, 44264, 44264, 44237, 44237, 44237, 44215, 44215, 44215, 44215, 44187, 44187, 44187, 44165, 44165, 44165, 44165, 44137, 44137, 44137, 44115, 44115, 44115, 44115, 44087, 44087, 44087, 44065, 44065, 44065, 44065, 44037, 44037, 44037, 44015, 44015, 44015, 44015, 43988, 43988, 43988, 43966, 43966, 43966, 43966, 43938, 43938, 43938, 43916, 43916, 43916, 43916, 43888, 43888, 43888, 43888, 43866, 43866, 43866, 43838, 43838, 43838, 43838, 43816, 43816, 43816, 43789, 43789, 43789, 43789, 43767, 43767, 43767, 43739, 43739, 43739, 43739, 43717, 43717, 43717, 43689, 43689, 43689, 43689, 43667, 43667, 43667, 43645, 43645, 43645, 43645, 43617, 43617, 43617, 43595, 43595, 43595, 43595, 43568, 43568, 43568, 43546, 43546, 43546, 43546, 43518, 43518, 43518, 43518, 43496, 43496, 43496, 43468, 43468, 43468, 43468, 43446, 43446, 43446, 43419, 43419, 43419, 43419, 43397, 43397, 43397, 43369, 43369, 43369, 43369, 43347, 43347, 43347, 43319, 43319, 43319, 43319, 43297, 43297, 43297, 43270, 43270, 43270, 43270, 43248, 43248, 43248, 43248, 43220, 43220, 43220, 43198, 43198, 43198, 43198, 43170, 43170, 43170, 43148, 43148, 43148, 43148, 43121, 43121, 43121, 43099, 43099, 43099, 43099, 43071, 43071, 43071, 43049, 43049, 43049, 43049, 43022, 43022, 43022, 43022, 43000, 43000, 43000, 42972, 42972, 42972, 42972, 42950, 42950, 42950, 42922, 42922, 42922, 42922, 42900, 42900, 42900, 42873, 42873, 42873, 42873, 42851, 42851, 42851, 42823, 42823, 42823, 42823, 42801, 42801, 42801, 42801, 42774, 42774, 42774, 42752, 42752, 42752, 42752, 42724, 42724, 42724, 42702, 42702, 42702, 42702, 42675, 42675, 42675, 42653, 42653, 42653, 42653, 42625, 42625, 42625, 42625, 42603, 42603, 42603, 42576, 42576, 42576, 42576, 42554, 42554, 42554, 42532, 42532, 42532, 42532, 42504, 42504, 42504, 42482, 42482, 42482, 42482, 42455, 42455, 42455, 42455, 42433, 42433, 42433, 42405, 42405, 42405, 42405, 42383, 42383, 42383, 42356, 42356, 42356, 42356, 42334, 42334, 42334, 42306, 42306, 42306, 42306, 42284, 42284, 42284, 42284, 42257, 42257, 42257, 42235, 42235, 42235, 42235, 42207, 42207, 42207, 42185, 42185, 42185, 42185, 42158, 42158, 42158, 42158, 42136, 42136, 42136, 42108, 42108, 42108, 42108, 42086, 42086, 42086, 42059, 42059, 42059, 42059, 42037, 42037, 42037, 42009, 42009, 42009, 42009, 41988, 41988, 41988, 41988, 41960, 41960, 41960, 41938, 41938, 41938, 41938, 41911, 41911, 41911, 41889, 41889, 41889, 41889, 41861, 41861, 41861, 41861, 41839, 41839, 41839, 41812, 41812, 41812, 41812, 41790, 41790, 41790, 41762, 41762, 41762, 41762, 41740, 41740, 41740, 41740, 41713, 41713, 41713, 41691, 41691, 41691, 41691, 41664, 41664, 41664, 41642, 41642, 41642, 41642, 41614, 41614, 41614, 41614, 41592, 41592, 41592, 41565, 41565, 41565, 41565, 41543, 41543, 41543, 41516, 41516, 41516, 41516, 41494, 41494, 41494, 41494, 41466, 41466, 41466, 41444, 41444, 41444, 41444, 41422, 41422, 41422, 41395, 41395, 41395, 41395, 41373, 41373, 41373, 41373, 41346, 41346, 41346, 41324, 41324, 41324, 41324, 41296, 41296, 41296, 41296, 41274, 41274, 41274, 41247, 41247, 41247, 41247, 41225, 41225, 41225, 41198, 41198, 41198, 41198, 41176, 41176, 41176, 41176, 41148, 41148, 41148, 41126, 41126, 41126, 41126, 41099, 41099, 41099, 41099, 41077, 41077, 41077, 41050, 41050, 41050, 41050, 41028, 41028, 41028, 41000, 41000, 41000, 41000, 40979, 40979, 40979, 40979, 40951, 40951, 40951, 40929, 40929, 40929, 40929, 40902, 40902, 40902, 40902, 40880, 40880, 40880, 40853, 40853, 40853, 40853, 40831, 40831, 40831, 40803, 40803, 40803, 40803, 40781, 40781, 40781, 40781, 40754, 40754, 40754, 40732, 40732, 40732, 40732, 40705, 40705, 40705, 40705, 40683, 40683, 40683, 40656, 40656, 40656, 40656, 40634, 40634, 40634, 40634, 40606, 40606, 40606, 40584, 40584, 40584, 40584, 40557, 40557, 40557, 40535, 40535, 40535, 40535, 40508, 40508, 40508, 40508, 40486, 40486, 40486, 40459, 40459, 40459, 40459, 40437, 40437, 40437, 40437, 40409, 40409, 40409, 40388, 40388, 40388, 40388, 40360, 40360, 40360, 40360, 40338, 40338, 40338, 40316, 40316, 40316, 40316, 40289, 40289, 40289, 40289, 40267, 40267, 40267, 40240, 40240, 40240, 40240, 40218, 40218, 40218, 40218, 40191, 40191, 40191, 40169, 40169, 40169, 40169, 40142, 40142, 40142, 40142, 40120, 40120, 40120, 40092, 40092, 40092, 40092, 40070, 40070, 40070, 40070, 40043, 40043, 40043, 40021, 40021, 40021, 40021, 39994, 39994, 39994, 39994, 39972, 39972, 39972, 39945, 39945, 39945, 39945, 39923, 39923, 39923, 39923, 39896, 39896, 39896, 39874, 39874, 39874, 39874, 39846, 39846, 39846, 39846, 39825, 39825, 39825, 39797, 39797, 39797, 39797, 39775, 39775, 39775, 39775, 39748, 39748, 39748, 39726, 39726, 39726, 39726, 39699, 39699, 39699, 39699, 39677, 39677, 39677, 39650, 39650, 39650, 39650, 39628, 39628, 39628, 39628, 39601, 39601, 39601, 39579, 39579, 39579, 39579, 39552, 39552, 39552, 39552, 39530, 39530, 39530, 39502, 39502, 39502, 39502, 39481, 39481, 39481, 39481, 39453, 39453, 39453, 39432, 39432, 39432, 39432, 39404, 39404, 39404, 39404, 39382, 39382, 39382, 39355, 39355, 39355, 39355, 39333, 39333, 39333, 39333, 39306, 39306, 39306, 39284, 39284, 39284, 39284, 39262, 39262, 39262, 39262, 39235, 39235, 39235, 39235, 39213, 39213, 39213, 39186, 39186, 39186, 39186, 39164, 39164, 39164, 39164, 39137, 39137, 39137, 39115, 39115, 39115, 39115, 39088, 39088, 39088, 39088, 39066, 39066, 39066, 39039, 39039, 39039, 39039, 39017, 39017, 39017, 39017, 38990, 38990, 38990, 38990, 38968, 38968, 38968, 38941, 38941, 38941, 38941, 38919, 38919, 38919, 38919, 38891, 38891, 38891, 38870, 38870, 38870, 38870, 38842, 38842, 38842, 38842, 38821, 38821, 38821, 38821, 38793, 38793, 38793, 38771, 38771, 38771, 38771, 38744, 38744, 38744, 38744, 38722, 38722, 38722, 38695, 38695, 38695, 38695, 38673, 38673, 38673, 38673, 38646, 38646, 38646, 38646, 38624, 38624, 38624, 38597, 38597, 38597, 38597, 38575, 38575, 38575, 38575, 38548, 38548, 38548, 38526, 38526, 38526, 38526, 38499, 38499, 38499, 38499, 38477, 38477, 38477, 38477, 38450, 38450, 38450, 38428, 38428, 38428, 38428, 38401, 38401, 38401, 38401, 38379, 38379, 38379, 38352, 38352, 38352, 38352, 38330, 38330, 38330, 38330, 38303, 38303, 38303, 38303, 38281, 38281, 38281, 38254, 38254, 38254, 38254, 38232, 38232, 38232, 38232, 38205, 38205, 38205, 38205, 38183, 38183, 38183, 38161, 38161, 38161, 38161, 38134, 38134, 38134, 38134, 38112, 38112, 38112, 38112, 38085, 38085, 38085, 38063, 38063, 38063, 38063, 38036, 38036, 38036, 38036, 38014, 38014, 38014, 38014, 37987, 37987, 37987, 37965, 37965, 37965, 37965, 37938, 37938, 37938, 37938, 37916, 37916, 37916, 37916, 37889, 37889, 37889, 37867, 37867, 37867, 37867, 37840, 37840, 37840, 37840, 37818, 37818, 37818, 37818, 37791, 37791, 37791, 37769, 37769, 37769, 37769, 37742, 37742, 37742, 37742, 37720, 37720, 37720, 37720, 37693, 37693, 37693, 37671, 37671, 37671, 37671, 37644, 37644, 37644, 37644, 37622, 37622, 37622, 37622, 37595, 37595, 37595, 37573, 37573, 37573, 37573, 37546, 37546, 37546, 37546, 37524, 37524, 37524, 37524, 37497, 37497, 37497, 37475, 37475, 37475, 37475, 37448, 37448, 37448, 37448, 37426, 37426, 37426, 37426, 37399, 37399, 37399, 37377, 37377, 37377, 37377, 37350, 37350, 37350, 37350, 37328, 37328, 37328, 37328, 37301, 37301, 37301, 37301, 37279, 37279, 37279, 37252, 37252, 37252, 37252, 37230, 37230, 37230, 37230, 37203, 37203, 37203, 37203, 37181, 37181, 37181, 37154, 37154, 37154, 37154, 37132, 37132, 37132, 37132, 37105, 37105, 37105, 37105, 37083, 37083, 37083, 37083, 37061, 37061, 37061, 37034, 37034, 37034, 37034, 37012, 37012, 37012, 37012, 36985, 36985, 36985, 36985, 36963, 36963, 36963, 36963, 36936, 36936, 36936, 36914, 36914, 36914, 36914, 36887, 36887, 36887, 36887, 36865, 36865, 36865, 36865, 36838, 36838, 36838, 36816, 36816, 36816, 36816, 36789, 36789, 36789, 36789, 36767, 36767, 36767, 36767, 36740, 36740, 36740, 36740, 36718, 36718, 36718, 36691, 36691, 36691, 36691, 36669, 36669, 36669, 36669, 36642, 36642, 36642, 36642, 36620, 36620, 36620, 36620, 36593, 36593, 36593, 36593, 36571, 36571, 36571, 36544, 36544, 36544, 36544, 36522, 36522, 36522, 36522, 36495, 36495, 36495, 36495, 36473, 36473, 36473, 36473, 36446, 36446, 36446, 36424, 36424, 36424, 36424, 36397, 36397, 36397, 36397, 36375, 36375, 36375, 36375, 36348, 36348, 36348, 36348, 36326, 36326, 36326, 36299, 36299, 36299, 36299, 36278, 36278, 36278, 36278, 36250, 36250, 36250, 36250, 36229, 36229, 36229, 36229, 36201, 36201, 36201, 36201, 36180, 36180, 36180, 36152, 36152, 36152, 36152, 36131, 36131, 36131, 36131, 36103, 36103, 36103, 36103, 36082, 36082, 36082, 36082, 36054, 36054, 36054, 36054, 36033, 36033, 36033, 36005, 36005, 36005, 36005, 35984, 35984, 35984, 35984, 35962, 35962, 35962, 35962, 35935, 35935, 35935, 35935, 35913, 35913, 35913, 35913, 35886, 35886, 35886, 35864, 35864, 35864, 35864, 35837, 35837, 35837, 35837, 35815, 35815, 35815, 35815, 35788, 35788, 35788, 35788, 35766, 35766, 35766, 35766, 35739, 35739, 35739, 35717, 35717, 35717, 35717, 35690, 35690, 35690, 35690, 35668, 35668, 35668, 35668, 35641, 35641, 35641, 35641, 35619, 35619, 35619, 35619, 35592, 35592, 35592, 35592, 35570, 35570, 35570, 35543, 35543, 35543, 35543, 35521, 35521, 35521, 35521, 35494, 35494, 35494, 35494, 35472, 35472, 35472, 35472, 35445, 35445, 35445, 35445, 35423, 35423, 35423, 35423, 35396, 35396, 35396, 35374, 35374, 35374, 35374, 35347, 35347, 35347, 35347, 35325, 35325, 35325, 35325, 35298, 35298, 35298, 35298, 35276, 35276, 35276, 35276, 35249, 35249, 35249, 35249, 35227, 35227, 35227, 35200, 35200, 35200, 35200, 35178, 35178, 35178, 35178, 35151, 35151, 35151, 35151, 35129, 35129, 35129, 35129, 35102, 35102, 35102, 35102, 35080, 35080, 35080, 35080, 35053, 35053, 35053, 35053, 35031, 35031, 35031, 35031, 35004, 35004, 35004, 34982, 34982, 34982, 34982, 34955, 34955, 34955, 34955, 34933, 34933, 34933, 34933, 34912, 34912, 34912, 34912, 34884, 34884, 34884, 34884, 34863, 34863, 34863, 34863, 34835, 34835, 34835, 34835, 34814, 34814, 34814, 34786, 34786, 34786, 34786, 34765, 34765, 34765, 34765, 34737, 34737, 34737, 34737, 34716, 34716, 34716, 34716, 34688, 34688, 34688, 34688, 34667, 34667, 34667, 34667, 34639, 34639, 34639, 34639, 34618, 34618, 34618, 34618, 34590, 34590, 34590, 34590, 34569, 34569, 34569, 34541, 34541, 34541, 34541, 34520, 34520, 34520, 34520, 34492, 34492, 34492, 34492, 34471, 34471, 34471, 34471, 34443, 34443, 34443, 34443, 34422, 34422, 34422, 34422, 34394, 34394, 34394, 34394, 34373, 34373, 34373, 34373, 34345, 34345, 34345, 34345, 34324, 34324, 34324, 34324, 34296, 34296, 34296, 34275, 34275, 34275, 34275, 34247, 34247, 34247, 34247, 34226, 34226, 34226, 34226, 34198, 34198, 34198, 34198, 34177, 34177, 34177, 34177, 34149, 34149, 34149, 34149, 34128, 34128, 34128, 34128, 34100, 34100, 34100, 34100, 34079, 34079, 34079, 34079, 34051, 34051, 34051, 34051, 34030, 34030, 34030, 34030, 34002, 34002, 34002, 34002, 33981, 33981, 33981, 33981, 33953, 33953, 33953, 33932, 33932, 33932, 33932, 33904, 33904, 33904, 33904, 33882, 33882, 33882, 33882, 33855, 33855, 33855, 33855, 33833, 33833, 33833, 33833, 33812, 33812, 33812, 33812, 33784, 33784, 33784, 33784, 33763, 33763, 33763, 33763, 33735, 33735, 33735, 33735, 33714, 33714, 33714, 33714, 33686, 33686, 33686, 33686, 33665, 33665, 33665, 33665, 33637, 33637, 33637, 33637, 33616, 33616, 33616, 33616, 33588, 33588, 33588, 33588, 33566, 33566, 33566, 33566, 33539, 33539, 33539, 33539, 33517, 33517, 33517, 33517, 33490, 33490, 33490, 33468, 33468, 33468, 33468, 33441, 33441, 33441, 33441, 33419, 33419, 33419, 33419, 33392, 33392, 33392, 33392, 33370, 33370, 33370, 33370, 33343, 33343, 33343, 33343, 33321, 33321, 33321, 33321, 33294, 33294, 33294, 33294, 33272, 33272, 33272, 33272, 33245, 33245, 33245, 33245, 33223, 33223, 33223, 33223, 33196, 33196, 33196, 33196, 33174, 33174, 33174, 33174, 33147, 33147, 33147, 33147, 33125, 33125, 33125, 33125, 33098, 33098, 33098, 33098, 33076, 33076, 33076, 33076, 33049, 33049, 33049, 33049, 33027, 33027, 33027, 33027, 32999, 32999, 32999, 32999, 32978, 32978, 32978, 32978, 32950, 32950, 32950, 32950, 32929, 32929, 32929, 32929, 32901, 32901, 32901, 32901, 32879, 32879, 32879, 32879, 32852, 32852, 32852, 32852, 32830, 32830, 32830, 32830, 32803, 32803, 32803, 32803, 32781, 32781, 32781, 32781, 32754, 32754, 32754, 32754, 32732, 32732, 32732, 32732, 32710, 32710, 32710, 32710, 32683, 32683, 32683, 32683, 32661, 32661, 32661, 32661, 32634, 32634, 32634, 32634, 32612, 32612, 32612, 32612, 32585, 32585, 32585, 32585, 32563, 32563, 32563, 32563, 32536, 32536, 32536, 32536, 32514, 32514, 32514, 32514, 32487, 32487, 32487, 32487, 32465, 32465, 32465, 32465, 32437, 32437, 32437, 32437, 32416, 32416, 32416, 32416, 32388, 32388, 32388, 32388, 32366, 32366, 32366, 32366, 32339, 32339, 32339, 32339, 32317, 32317, 32317, 32317, 32290, 32290, 32290, 32290, 32268, 32268, 32268, 32268, 32241, 32241, 32241, 32241, 32219, 32219, 32219, 32219, 32192, 32192, 32192, 32192, 32170, 32170, 32170, 32170, 32143, 32143, 32143, 32143, 32121, 32121, 32121, 32121, 32093, 32093, 32093, 32093, 32072, 32072, 32072, 32072, 32044, 32044, 32044, 32044, 32044, 32022, 32022, 32022, 32022, 31995, 31995, 31995, 31995, 31973, 31973, 31973, 31973, 31946, 31946, 31946, 31946, 31924, 31924, 31924, 31924, 31897, 31897, 31897, 31897, 31875, 31875, 31875, 31875, 31848, 31848, 31848, 31848, 31826, 31826, 31826, 31826, 31798, 31798, 31798, 31798, 31776, 31776, 31776, 31776, 31749, 31749, 31749, 31749, 31727, 31727, 31727, 31727, 31700, 31700, 31700, 31700, 31678, 31678, 31678, 31678, 31651, 31651, 31651, 31651, 31629, 31629, 31629, 31629, 31607, 31607, 31607, 31607, 31580, 31580, 31580, 31580, 31580, 31558, 31558, 31558, 31558, 31530, 31530, 31530, 31530, 31509, 31509, 31509, 31509, 31481, 31481, 31481, 31481, 31459, 31459, 31459, 31459, 31432, 31432, 31432, 31432, 31410, 31410, 31410, 31410, 31383, 31383, 31383, 31383, 31361, 31361, 31361, 31361, 31333, 31333, 31333, 31333, 31312, 31312, 31312, 31312, 31284, 31284, 31284, 31284, 31262, 31262, 31262, 31262, 31262, 31235, 31235, 31235, 31235, 31213, 31213, 31213, 31213, 31186, 31186, 31186, 31186, 31164, 31164, 31164, 31164, 31136, 31136, 31136, 31136, 31115, 31115, 31115, 31115, 31087, 31087, 31087, 31087, 31065, 31065, 31065, 31065, 31038, 31038, 31038, 31038, 31016, 31016, 31016, 31016, 31016, 30989, 30989, 30989, 30989, 30967, 30967, 30967, 30967, 30939, 30939, 30939, 30939, 30917, 30917, 30917, 30917, 30890, 30890, 30890, 30890, 30868, 30868, 30868, 30868, 30841, 30841, 30841, 30841, 30819, 30819, 30819, 30819, 30791, 30791, 30791, 30791, 30791, 30769, 30769, 30769, 30769, 30742, 30742, 30742, 30742, 30720, 30720, 30720, 30720, 30693, 30693, 30693, 30693, 30671, 30671, 30671, 30671, 30643, 30643, 30643, 30643, 30622, 30622, 30622, 30622, 30594, 30594, 30594, 30594, 30572, 30572, 30572, 30572, 30572, 30545, 30545, 30545, 30545, 30523, 30523, 30523, 30523, 30501, 30501, 30501, 30501, 30473, 30473, 30473, 30473, 30452, 30452, 30452, 30452, 30424, 30424, 30424, 30424, 30402, 30402, 30402, 30402, 30402, 30375, 30375, 30375, 30375, 30353, 30353, 30353, 30353, 30325, 30325, 30325, 30325, 30303, 30303, 30303, 30303, 30276, 30276, 30276, 30276, 30254, 30254, 30254, 30254, 30227, 30227, 30227, 30227, 30227, 30205, 30205, 30205, 30205, 30177, 30177, 30177, 30177, 30155, 30155, 30155, 30155, 30128, 30128, 30128, 30128, 30106, 30106, 30106, 30106, 30078, 30078, 30078, 30078, 30078, 30056, 30056, 30056, 30056, 30029, 30029, 30029, 30029, 30007, 30007, 30007, 30007, 29980, 29980, 29980, 29980, 29958, 29958, 29958, 29958, 29930, 29930, 29930, 29930, 29930, 29908, 29908, 29908, 29908, 29881, 29881, 29881, 29881, 29859, 29859, 29859, 29859, 29831, 29831, 29831, 29831, 29809, 29809, 29809, 29809, 29782, 29782, 29782, 29782, 29782, 29760, 29760, 29760, 29760, 29732, 29732, 29732, 29732, 29710, 29710, 29710, 29710, 29683, 29683, 29683, 29683, 29661, 29661, 29661, 29661, 29661, 29633, 29633, 29633, 29633, 29611, 29611, 29611, 29611, 29584, 29584, 29584, 29584, 29562, 29562, 29562, 29562, 29534, 29534, 29534, 29534, 29534, 29512, 29512, 29512, 29512, 29485, 29485, 29485, 29485, 29463, 29463, 29463, 29463, 29441, 29441, 29441, 29441, 29413, 29413, 29413, 29413, 29413, 29391, 29391, 29391, 29391, 29364, 29364, 29364, 29364, 29342, 29342, 29342, 29342, 29314, 29314, 29314, 29314, 29292, 29292, 29292, 29292, 29292, 29265, 29265, 29265, 29265, 29243, 29243, 29243, 29243, 29215, 29215, 29215, 29215, 29193, 29193, 29193, 29193, 29166, 29166, 29166, 29166, 29166, 29144, 29144, 29144, 29144, 29116, 29116, 29116, 29116, 29094, 29094, 29094, 29094, 29066, 29066, 29066, 29066, 29066, 29044, 29044, 29044, 29044, 29017, 29017, 29017, 29017, 28995, 28995, 28995, 28995, 28967, 28967, 28967, 28967, 28967, 28945, 28945, 28945, 28945, 28918, 28918, 28918, 28918, 28896, 28896, 28896, 28896, 28868, 28868, 28868, 28868, 28846, 28846, 28846, 28846, 28846, 28818, 28818, 28818, 28818, 28796, 28796, 28796, 28796, 28769, 28769, 28769, 28769, 28747, 28747, 28747, 28747, 28747, 28719, 28719, 28719, 28719, 28697, 28697, 28697, 28697, 28670, 28670, 28670, 28670, 28648, 28648, 28648, 28648, 28648, 28620, 28620, 28620, 28620, 28598, 28598, 28598, 28598, 28570, 28570, 28570, 28570, 28570, 28548, 28548, 28548, 28548, 28521, 28521, 28521, 28521, 28499, 28499, 28499, 28499, 28471, 28471, 28471, 28471, 28471, 28449, 28449, 28449, 28449, 28421, 28421, 28421, 28421, 28399, 28399, 28399, 28399, 28372, 28372, 28372, 28372, 28372, 28349, 28349, 28349, 28349, 28327, 28327, 28327, 28327, 28300, 28300, 28300, 28300, 28300, 28278, 28278, 28278, 28278, 28250, 28250, 28250, 28250, 28228, 28228, 28228, 28228, 28200, 28200, 28200, 28200, 28200, 28178, 28178, 28178, 28178, 28151, 28151, 28151, 28151, 28128, 28128, 28128, 28128, 28128, 28101, 28101, 28101, 28101, 28079, 28079, 28079, 28079, 28051, 28051, 28051, 28051, 28029, 28029, 28029, 28029, 28029, 28001, 28001, 28001, 28001, 27979, 27979, 27979, 27979, 27951, 27951, 27951, 27951, 27951, 27929, 27929, 27929, 27929, 27902, 27902, 27902, 27902, 27880, 27880, 27880, 27880, 27880, 27852, 27852, 27852, 27852, 27830, 27830, 27830, 27830, 27802, 27802, 27802, 27802, 27802, 27780, 27780, 27780, 27780, 27752, 27752, 27752, 27752, 27730, 27730, 27730, 27730, 27730, 27702, 27702, 27702, 27702, 27680, 27680, 27680, 27680, 27653, 27653, 27653, 27653, 27653, 27630, 27630, 27630, 27630, 27603, 27603, 27603, 27603, 27581, 27581, 27581, 27581, 27581, 27553, 27553, 27553, 27553, 27531, 27531, 27531, 27531, 27503, 27503, 27503, 27503, 27503, 27481, 27481, 27481, 27481, 27453, 27453, 27453, 27453, 27431, 27431, 27431, 27431, 27431, 27403, 27403, 27403, 27403, 27381, 27381, 27381, 27381, 27353, 27353, 27353, 27353, 27353, 27331, 27331, 27331, 27331, 27303, 27303, 27303, 27303, 27281, 27281, 27281, 27281, 27281, 27253, 27253, 27253, 27253, 27231, 27231, 27231, 27231, 27209, 27209, 27209, 27209, 27209, 27181, 27181, 27181, 27181, 27159, 27159, 27159, 27159, 27159, 27131, 27131, 27131, 27131, 27109, 27109, 27109, 27109, 27081, 27081, 27081, 27081, 27081, 27059, 27059, 27059, 27059, 27031, 27031, 27031, 27031, 27009, 27009, 27009, 27009, 27009, 26981, 26981, 26981, 26981, 26959, 26959, 26959, 26959, 26959, 26931, 26931, 26931, 26931, 26909, 26909, 26909, 26909, 26881, 26881, 26881, 26881, 26881, 26859, 26859, 26859, 26859, 26831, 26831, 26831, 26831, 26831, 26809, 26809, 26809, 26809, 26781, 26781, 26781, 26781, 26759, 26759, 26759, 26759, 26759, 26731, 26731, 26731, 26731, 26709, 26709, 26709, 26709, 26709, 26681, 26681, 26681, 26681, 26659, 26659, 26659, 26659, 26631, 26631, 26631, 26631, 26631, 26609, 26609, 26609, 26609, 26581, 26581, 26581, 26581, 26581, 26559, 26559, 26559, 26559, 26531, 26531, 26531, 26531, 26509, 26509, 26509, 26509, 26509, 26481, 26481, 26481, 26481, 26459, 26459, 26459, 26459, 26459, 26431, 26431, 26431, 26431, 26408, 26408, 26408, 26408, 26408, 26381, 26381, 26381, 26381, 26358, 26358, 26358, 26358, 26330, 26330, 26330, 26330, 26330, 26308, 26308, 26308, 26308, 26280, 26280, 26280, 26280, 26280, 26258, 26258, 26258, 26258, 26230, 26230, 26230, 26230, 26230, 26208, 26208, 26208, 26208, 26180, 26180, 26180, 26180, 26158, 26158, 26158, 26158, 26158, 26130, 26130, 26130, 26130, 26107, 26107, 26107, 26107, 26107, 26085, 26085, 26085, 26085, 26057, 26057, 26057, 26057, 26057, 26035, 26035, 26035, 26035, 26007, 26007, 26007, 26007, 26007, 25985, 25985, 25985, 25985, 25957, 25957, 25957, 25957, 25957, 25934, 25934, 25934, 25934, 25906, 25906, 25906, 25906, 25884, 25884, 25884, 25884, 25884, 25856, 25856, 25856, 25856, 25834, 25834, 25834, 25834, 25834, 25806, 25806, 25806, 25806, 25784, 25784, 25784, 25784, 25784, 25756, 25756, 25756, 25756, 25733, 25733, 25733, 25733, 25733, 25705, 25705, 25705, 25705, 25683, 25683, 25683, 25683, 25683, 25655, 25655, 25655, 25655, 25633, 25633, 25633, 25633, 25633, 25605, 25605, 25605, 25605, 25582, 25582, 25582, 25582, 25582, 25554, 25554, 25554, 25554, 25532, 25532, 25532, 25532, 25532, 25504, 25504, 25504, 25504, 25482, 25482, 25482, 25482, 25482, 25454, 25454, 25454, 25454, 25431, 25431, 25431, 25431, 25431, 25403, 25403, 25403, 25403, 25381, 25381, 25381, 25381, 25381, 25353, 25353, 25353, 25353, 25330, 25330, 25330, 25330, 25330, 25302, 25302, 25302, 25302, 25280, 25280, 25280, 25280, 25280, 25252, 25252, 25252, 25252, 25230, 25230, 25230, 25230, 25230, 25202, 25202, 25202, 25202, 25179, 25179, 25179, 25179, 25179, 25151, 25151, 25151, 25151, 25151, 25129, 25129, 25129, 25129, 25101, 25101, 25101, 25101, 25101, 25078, 25078, 25078, 25078, 25050, 25050, 25050, 25050, 25050, 25028, 25028, 25028, 25028, 25005, 25005, 25005, 25005, 25005, 24977, 24977, 24977, 24977, 24955, 24955, 24955, 24955, 24955, 24927, 24927, 24927, 24927, 24904, 24904, 24904, 24904, 24904, 24876, 24876, 24876, 24876, 24876, 24854, 24854, 24854, 24854, 24826, 24826, 24826, 24826, 24826, 24803, 24803, 24803, 24803, 24775, 24775, 24775, 24775, 24775, 24753, 24753, 24753, 24753, 24725, 24725, 24725, 24725, 24725, 24702, 24702, 24702, 24702, 24702, 24674, 24674, 24674, 24674, 24652, 24652, 24652, 24652, 24652, 24623, 24623, 24623, 24623, 24601, 24601, 24601, 24601, 24601, 24573, 24573, 24573, 24573, 24550, 24550, 24550, 24550, 24550, 24522, 24522, 24522, 24522, 24522, 24500, 24500, 24500, 24500, 24472, 24472, 24472, 24472, 24472, 24449, 24449, 24449, 24449, 24421, 24421, 24421, 24421, 24421, 24398, 24398, 24398, 24398, 24398, 24370, 24370, 24370, 24370, 24348, 24348, 24348, 24348, 24348, 24320, 24320, 24320, 24320, 24297, 24297, 24297, 24297, 24297, 24269, 24269, 24269, 24269, 24269, 24246, 24246, 24246, 24246, 24218, 24218, 24218, 24218, 24218, 24196, 24196, 24196, 24196, 24167, 24167, 24167, 24167, 24167, 24145, 24145, 24145, 24145, 24145, 24117, 24117, 24117, 24117, 24094, 24094, 24094, 24094, 24094, 24066, 24066, 24066, 24066, 24066, 24043, 24043, 24043, 24043, 24015, 24015, 24015, 24015, 24015, 23993, 23993, 23993, 23993, 23993, 23964, 23964, 23964, 23964, 23942, 23942, 23942, 23942, 23942, 23914, 23914, 23914, 23914, 23891, 23891, 23891, 23891, 23891, 23868, 23868, 23868, 23868, 23868, 23840, 23840, 23840, 23840, 23818, 23818, 23818, 23818, 23818, 23789, 23789, 23789, 23789, 23789, 23767, 23767, 23767, 23767, 23738, 23738, 23738, 23738, 23738, 23716, 23716, 23716, 23716, 23716, 23688, 23688, 23688, 23688, 23665, 23665, 23665, 23665, 23665, 23637, 23637, 23637, 23637, 23637, 23614, 23614, 23614, 23614, 23586, 23586, 23586, 23586, 23586, 23563, 23563, 23563, 23563, 23563, 23535, 23535, 23535, 23535, 23512, 23512, 23512, 23512, 23512, 23484, 23484, 23484, 23484, 23484, 23461, 23461, 23461, 23461, 23461, 23433, 23433, 23433, 23433, 23410, 23410, 23410, 23410, 23410, 23382, 23382, 23382, 23382, 23382, 23359, 23359, 23359, 23359, 23331, 23331, 23331, 23331, 23331, 23308, 23308, 23308, 23308, 23308, 23280, 23280, 23280, 23280, 23257, 23257, 23257, 23257, 23257, 23229, 23229, 23229, 23229, 23229, 23206, 23206, 23206, 23206, 23206, 23178, 23178, 23178, 23178, 23155, 23155, 23155, 23155, 23155, 23127, 23127, 23127, 23127, 23127, 23104, 23104, 23104, 23104, 23076, 23076, 23076, 23076, 23076, 23053, 23053, 23053, 23053, 23053, 23025, 23025, 23025, 23025, 23025, 23002, 23002, 23002, 23002, 22974, 22974, 22974, 22974, 22974, 22951, 22951, 22951, 22951, 22951, 22922, 22922, 22922, 22922, 22922, 22900, 22900, 22900, 22900, 22871, 22871, 22871, 22871, 22871, 22849, 22849, 22849, 22849, 22849, 22820, 22820, 22820, 22820, 22820, 22797, 22797, 22797, 22797, 22769, 22769, 22769, 22769, 22769, 22746, 22746, 22746, 22746, 22746, 22724, 22724, 22724, 22724, 22724, 22695, 22695, 22695, 22695, 22672, 22672, 22672, 22672, 22672, 22644, 22644, 22644, 22644, 22644, 22621, 22621, 22621, 22621, 22621, 22593, 22593, 22593, 22593, 22593, 22570, 22570, 22570, 22570, 22541, 22541, 22541, 22541, 22541, 22519, 22519, 22519, 22519, 22519, 22490, 22490, 22490, 22490, 22490, 22467, 22467, 22467, 22467, 22439, 22439, 22439, 22439, 22439, 22416, 22416, 22416, 22416, 22416, 22388, 22388, 22388, 22388, 22388, 22365, 22365, 22365, 22365, 22365, 22336, 22336, 22336, 22336, 22313, 22313, 22313, 22313, 22313, 22285, 22285, 22285, 22285, 22285, 22262, 22262, 22262, 22262, 22262, 22234, 22234, 22234, 22234, 22234, 22211, 22211, 22211, 22211, 22211, 22182, 22182, 22182, 22182, 22159, 22159, 22159, 22159, 22159, 22131, 22131, 22131, 22131, 22131, 22108, 22108, 22108, 22108, 22108, 22079, 22079, 22079, 22079, 22079, 22057, 22057, 22057, 22057, 22057, 22028, 22028, 22028, 22028, 22005, 22005, 22005, 22005, 22005, 21977, 21977, 21977, 21977, 21977, 21954, 21954, 21954, 21954, 21954, 21925, 21925, 21925, 21925, 21925, 21902, 21902, 21902, 21902, 21902, 21874, 21874, 21874, 21874, 21851, 21851, 21851, 21851, 21851, 21822, 21822, 21822, 21822, 21822, 21799, 21799, 21799, 21799, 21799, 21771, 21771, 21771, 21771, 21771, 21748, 21748, 21748, 21748, 21748, 21719, 21719, 21719, 21719, 21719, 21696, 21696, 21696, 21696, 21696, 21668, 21668, 21668, 21668, 21645, 21645, 21645, 21645, 21645, 21616, 21616, 21616, 21616, 21616, 21593, 21593, 21593, 21593, 21593, 21570, 21570, 21570, 21570, 21570, 21541, 21541, 21541, 21541, 21541, 21518, 21518, 21518, 21518, 21518, 21490, 21490, 21490, 21490, 21490, 21467, 21467, 21467, 21467, 21467, 21438, 21438, 21438, 21438, 21415, 21415, 21415, 21415, 21415, 21387, 21387, 21387, 21387, 21387, 21364, 21364, 21364, 21364, 21364, 21335, 21335, 21335, 21335, 21335, 21312, 21312, 21312, 21312, 21312, 21283, 21283, 21283, 21283, 21283, 21260, 21260, 21260, 21260, 21260, 21231, 21231, 21231, 21231, 21231, 21208, 21208, 21208, 21208, 21208, 21180, 21180, 21180, 21180, 21180, 21157, 21157, 21157, 21157, 21157, 21128, 21128, 21128, 21128, 21128, 21105, 21105, 21105, 21105, 21076, 21076, 21076, 21076, 21076, 21053, 21053, 21053, 21053, 21053, 21024, 21024, 21024, 21024, 21024, 21001, 21001, 21001, 21001, 21001, 20973, 20973, 20973, 20973, 20973, 20950, 20950, 20950, 20950, 20950, 20921, 20921, 20921, 20921, 20921, 20898, 20898, 20898, 20898, 20898, 20869, 20869, 20869, 20869, 20869, 20846, 20846, 20846, 20846, 20846, 20817, 20817, 20817, 20817, 20817, 20794, 20794, 20794, 20794, 20794, 20765, 20765, 20765, 20765, 20765, 20742, 20742, 20742, 20742, 20742, 20713, 20713, 20713, 20713, 20713, 20690, 20690, 20690, 20690, 20690, 20661, 20661, 20661, 20661, 20661, 20638, 20638, 20638, 20638, 20638, 20609, 20609, 20609, 20609, 20609, 20586, 20586, 20586, 20586, 20586, 20557, 20557, 20557, 20557, 20557, 20534, 20534, 20534, 20534, 20534, 20505, 20505, 20505, 20505, 20505, 20482, 20482, 20482, 20482, 20482, 20453, 20453, 20453, 20453, 20453, 20430, 20430, 20430, 20430, 20430, 20407, 20407, 20407, 20407, 20407, 20378, 20378, 20378, 20378, 20378, 20355, 20355, 20355, 20355, 20355, 20326, 20326, 20326, 20326, 20326, 20303, 20303, 20303, 20303, 20303, 20274, 20274, 20274, 20274, 20274, 20251, 20251, 20251, 20251, 20251, 20222, 20222, 20222, 20222, 20222, 20199, 20199, 20199, 20199, 20199, 20170, 20170, 20170, 20170, 20170, 20147, 20147, 20147, 20147, 20147, 20147, 20118, 20118, 20118, 20118, 20118, 20095, 20095, 20095, 20095, 20095, 20066, 20066, 20066, 20066, 20066, 20042, 20042, 20042, 20042, 20042, 20013, 20013, 20013, 20013, 20013, 19990, 19990, 19990, 19990, 19990, 19961, 19961, 19961, 19961, 19961, 19938, 19938, 19938, 19938, 19938, 19909, 19909, 19909, 19909, 19909, 19886, 19886, 19886, 19886, 19886, 19857, 19857, 19857, 19857, 19857, 19834, 19834, 19834, 19834, 19834, 19805, 19805, 19805, 19805, 19805, 19805, 19781, 19781, 19781, 19781, 19781, 19752, 19752, 19752, 19752, 19752, 19729, 19729, 19729, 19729, 19729, 19700, 19700, 19700, 19700, 19700, 19677, 19677, 19677, 19677, 19677, 19648, 19648, 19648, 19648, 19648, 19624, 19624, 19624, 19624, 19624, 19595, 19595, 19595, 19595, 19595, 19595, 19572, 19572, 19572, 19572, 19572, 19543, 19543, 19543, 19543, 19543, 19520, 19520, 19520, 19520, 19520, 19490, 19490, 19490, 19490, 19490, 19467, 19467, 19467, 19467, 19467, 19438, 19438, 19438, 19438, 19438, 19415, 19415, 19415, 19415, 19415, 19415, 19386, 19386, 19386, 19386, 19386, 19362, 19362, 19362, 19362, 19362, 19333, 19333, 19333, 19333, 19333, 19310, 19310, 19310, 19310, 19310, 19287, 19287, 19287, 19287, 19287, 19257, 19257, 19257, 19257, 19257, 19257, 19234, 19234, 19234, 19234, 19234, 19205, 19205, 19205, 19205, 19205, 19181, 19181, 19181, 19181, 19181, 19152, 19152, 19152, 19152, 19152, 19129, 19129, 19129, 19129, 19129, 19100, 19100, 19100, 19100, 19100, 19100, 19076, 19076, 19076, 19076, 19076, 19047, 19047, 19047, 19047, 19047, 19024, 19024, 19024, 19024, 19024, 18995, 18995, 18995, 18995, 18995, 18971, 18971, 18971, 18971, 18971, 18971, 18942, 18942, 18942, 18942, 18942, 18919, 18919, 18919, 18919, 18919, 18889, 18889, 18889, 18889, 18889, 18866, 18866, 18866, 18866, 18866, 18866, 18837, 18837, 18837, 18837, 18837, 18813, 18813, 18813, 18813, 18813, 18784, 18784, 18784, 18784, 18784, 18760, 18760, 18760, 18760, 18760, 18760, 18731, 18731, 18731, 18731, 18731, 18708, 18708, 18708, 18708, 18708, 18678, 18678, 18678, 18678, 18678, 18655, 18655, 18655, 18655, 18655, 18655, 18626, 18626, 18626, 18626, 18626, 18602, 18602, 18602, 18602, 18602, 18573, 18573, 18573, 18573, 18573, 18549, 18549, 18549, 18549, 18549, 18549, 18520, 18520, 18520, 18520, 18520, 18497, 18497, 18497, 18497, 18497, 18467, 18467, 18467, 18467, 18467, 18444, 18444, 18444, 18444, 18444, 18444, 18414, 18414, 18414, 18414, 18414, 18391, 18391, 18391, 18391, 18391, 18362, 18362, 18362, 18362, 18362, 18362, 18338, 18338, 18338, 18338, 18338, 18309, 18309, 18309, 18309, 18309, 18285, 18285, 18285, 18285, 18285, 18285, 18256, 18256, 18256, 18256, 18256, 18232, 18232, 18232, 18232, 18232, 18203, 18203, 18203, 18203, 18203, 18179, 18179, 18179, 18179, 18179, 18179, 18150, 18150, 18150, 18150, 18150, 18126, 18126, 18126, 18126, 18126, 18103, 18103, 18103, 18103, 18103, 18103, 18073, 18073, 18073, 18073, 18073, 18050, 18050, 18050, 18050, 18050, 18050, 18020, 18020, 18020, 18020, 18020, 17997, 17997, 17997, 17997, 17997, 17967, 17967, 17967, 17967, 17967, 17967, 17944, 17944, 17944, 17944, 17944, 17914, 17914, 17914, 17914, 17914, 17890, 17890, 17890, 17890, 17890, 17890, 17861, 17861, 17861, 17861, 17861, 17837, 17837, 17837, 17837, 17837, 17808, 17808, 17808, 17808, 17808, 17808, 17784, 17784, 17784, 17784, 17784, 17755, 17755, 17755, 17755, 17755, 17755, 17731, 17731, 17731, 17731, 17731, 17701, 17701, 17701, 17701, 17701, 17678, 17678, 17678, 17678, 17678, 17678, 17648, 17648, 17648, 17648, 17648, 17625, 17625, 17625, 17625, 17625, 17625, 17595, 17595, 17595, 17595, 17595, 17571, 17571, 17571, 17571, 17571, 17542, 17542, 17542, 17542, 17542, 17542, 17518, 17518, 17518, 17518, 17518, 17489, 17489, 17489, 17489, 17489, 17489, 17465, 17465, 17465, 17465, 17465, 17435, 17435, 17435, 17435, 17435, 17435, 17412, 17412, 17412, 17412, 17412, 17382, 17382, 17382, 17382, 17382, 17358, 17358, 17358, 17358, 17358, 17358, 17329, 17329, 17329, 17329, 17329, 17305, 17305, 17305, 17305, 17305, 17305, 17275, 17275, 17275, 17275, 17275, 17251, 17251, 17251, 17251, 17251, 17251, 17222, 17222, 17222, 17222, 17222, 17198, 17198, 17198, 17198, 17198, 17198, 17168, 17168, 17168, 17168, 17168, 17145, 17145, 17145, 17145, 17145, 17145, 17115, 17115, 17115, 17115, 17115, 17091, 17091, 17091, 17091, 17091, 17091, 17061, 17061, 17061, 17061, 17061, 17038, 17038, 17038, 17038, 17038, 17038, 17008, 17008, 17008, 17008, 17008, 16984, 16984, 16984, 16984, 16984, 16984, 16954, 16954, 16954, 16954, 16954, 16931, 16931, 16931, 16931, 16931, 16931, 16907, 16907, 16907, 16907, 16907, 16877, 16877, 16877, 16877, 16877, 16877, 16853, 16853, 16853, 16853, 16853, 16823, 16823, 16823, 16823, 16823, 16823, 16800, 16800, 16800, 16800, 16800, 16770, 16770, 16770, 16770, 16770, 16770, 16746, 16746, 16746, 16746, 16746, 16716, 16716, 16716, 16716, 16716, 16716, 16692, 16692, 16692, 16692, 16692, 16692, 16662, 16662, 16662, 16662, 16662, 16639, 16639, 16639, 16639, 16639, 16639, 16609, 16609, 16609, 16609, 16609, 16585, 16585, 16585, 16585, 16585, 16585, 16555, 16555, 16555, 16555, 16555, 16531, 16531, 16531, 16531, 16531, 16531, 16501, 16501, 16501, 16501, 16501, 16501, 16477, 16477, 16477, 16477, 16477, 16448, 16448, 16448, 16448, 16448, 16448, 16424, 16424, 16424, 16424, 16424, 16394, 16394, 16394, 16394, 16394, 16394, 16370, 16370, 16370, 16370, 16370, 16370, 16340, 16340, 16340, 16340, 16340, 16316, 16316, 16316, 16316, 16316, 16316, 16286, 16286, 16286, 16286, 16286, 16286, 16262, 16262, 16262, 16262, 16262, 16232, 16232, 16232, 16232, 16232, 16232, 16208, 16208, 16208, 16208, 16208, 16178, 16178, 16178, 16178, 16178, 16178, 16154, 16154, 16154, 16154, 16154, 16154, 16124, 16124, 16124, 16124, 16124, 16100, 16100, 16100, 16100, 16100, 16100, 16070, 16070, 16070, 16070, 16070, 16070, 16046, 16046, 16046, 16046, 16046, 16016, 16016, 16016, 16016, 16016, 16016, 15992, 15992, 15992, 15992, 15992, 15992, 15962, 15962, 15962, 15962, 15962, 15938, 15938, 15938, 15938, 15938, 15938, 15908, 15908, 15908, 15908, 15908, 15908, 15884, 15884, 15884, 15884, 15884, 15884, 15854, 15854, 15854, 15854, 15854, 15830, 15830, 15830, 15830, 15830, 15830, 15800, 15800, 15800, 15800, 15800, 15800, 15776, 15776, 15776, 15776, 15776, 15746, 15746, 15746, 15746, 15746, 15746, 15722, 15722, 15722, 15722, 15722, 15722, 15698, 15698, 15698, 15698, 15698, 15698, 15668, 15668, 15668, 15668, 15668, 15644, 15644, 15644, 15644, 15644, 15644, 15614, 15614, 15614, 15614, 15614, 15614, 15590, 15590, 15590, 15590, 15590, 15590, 15559, 15559, 15559, 15559, 15559, 15535, 15535, 15535, 15535, 15535, 15535, 15505, 15505, 15505, 15505, 15505, 15505, 15481, 15481, 15481, 15481, 15481, 15481, 15451, 15451, 15451, 15451, 15451, 15427, 15427, 15427, 15427, 15427, 15427, 15397, 15397, 15397, 15397, 15397, 15397, 15372, 15372, 15372, 15372, 15372, 15372, 15342, 15342, 15342, 15342, 15342, 15342, 15318, 15318, 15318, 15318, 15318, 15288, 15288, 15288, 15288, 15288, 15288, 15264, 15264, 15264, 15264, 15264, 15264, 15233, 15233, 15233, 15233, 15233, 15233, 15209, 15209, 15209, 15209, 15209, 15209, 15179, 15179, 15179, 15179, 15179, 15179, 15155, 15155, 15155, 15155, 15155, 15125, 15125, 15125, 15125, 15125, 15125, 15100, 15100, 15100, 15100, 15100, 15100, 15070, 15070, 15070, 15070, 15070, 15070, 15046, 15046, 15046, 15046, 15046, 15046, 15016, 15016, 15016, 15016, 15016, 15016, 14991, 14991, 14991, 14991, 14991, 14991, 14961, 14961, 14961, 14961, 14961, 14937, 14937, 14937, 14937, 14937, 14937, 14907, 14907, 14907, 14907, 14907, 14907, 14882, 14882, 14882, 14882, 14882, 14882, 14852, 14852, 14852, 14852, 14852, 14852, 14828, 14828, 14828, 14828, 14828, 14828, 14797, 14797, 14797, 14797, 14797, 14797, 14773, 14773, 14773, 14773, 14773, 14773, 14743, 14743, 14743, 14743, 14743, 14743, 14718, 14718, 14718, 14718, 14718, 14718, 14688, 14688, 14688, 14688, 14688, 14688, 14664, 14664, 14664, 14664, 14664, 14633, 14633, 14633, 14633, 14633, 14633, 14609, 14609, 14609, 14609, 14609, 14609, 14579, 14579, 14579, 14579, 14579, 14579, 14554, 14554, 14554, 14554, 14554, 14554, 14530, 14530, 14530, 14530, 14530, 14530, 14499, 14499, 14499, 14499, 14499, 14499, 14475, 14475, 14475, 14475, 14475, 14475, 14445, 14445, 14445, 14445, 14445, 14445, 14420, 14420, 14420, 14420, 14420, 14420, 14390, 14390, 14390, 14390, 14390, 14390, 14365, 14365, 14365, 14365, 14365, 14365, 14335, 14335, 14335, 14335, 14335, 14335, 14311, 14311, 14311, 14311, 14311, 14311, 14280, 14280, 14280, 14280, 14280, 14280, 14256, 14256, 14256, 14256, 14256, 14256, 14225, 14225, 14225, 14225, 14225, 14225, 14201, 14201, 14201, 14201, 14201, 14201, 14170, 14170, 14170, 14170, 14170, 14170, 14146, 14146, 14146, 14146, 14146, 14146, 14115, 14115, 14115, 14115, 14115, 14115, 14091, 14091, 14091, 14091, 14091, 14091, 14060, 14060, 14060, 14060, 14060, 14060, 14060, 14036, 14036, 14036, 14036, 14036, 14036, 14005, 14005, 14005, 14005, 14005, 14005, 13981, 13981, 13981, 13981, 13981, 13981, 13950, 13950, 13950, 13950, 13950, 13950, 13925, 13925, 13925, 13925, 13925, 13925, 13895, 13895, 13895, 13895, 13895, 13895, 13870, 13870, 13870, 13870, 13870, 13870, 13840, 13840, 13840, 13840, 13840, 13840, 13815, 13815, 13815, 13815, 13815, 13815, 13785, 13785, 13785, 13785, 13785, 13785, 13785, 13760, 13760, 13760, 13760, 13760, 13760, 13729, 13729, 13729, 13729, 13729, 13729, 13705, 13705, 13705, 13705, 13705, 13705, 13674, 13674, 13674, 13674, 13674, 13674, 13650, 13650, 13650, 13650, 13650, 13650, 13619, 13619, 13619, 13619, 13619, 13619, 13594, 13594, 13594, 13594, 13594, 13594, 13594, 13564, 13564, 13564, 13564, 13564, 13564, 13539, 13539, 13539, 13539, 13539, 13539, 13508, 13508, 13508, 13508, 13508, 13508, 13484, 13484, 13484, 13484, 13484, 13484, 13453, 13453, 13453, 13453, 13453, 13453, 13453, 13428, 13428, 13428, 13428, 13428, 13428, 13397, 13397, 13397, 13397, 13397, 13397, 13373, 13373, 13373, 13373, 13373, 13373, 13342, 13342, 13342, 13342, 13342, 13342, 13317, 13317, 13317, 13317, 13317, 13317, 13317, 13293, 13293, 13293, 13293, 13293, 13293, 13262, 13262, 13262, 13262, 13262, 13262, 13237, 13237, 13237, 13237, 13237, 13237, 13206, 13206, 13206, 13206, 13206, 13206, 13206, 13182, 13182, 13182, 13182, 13182, 13182, 13151, 13151, 13151, 13151, 13151, 13151, 13126, 13126, 13126, 13126, 13126, 13126, 13095, 13095, 13095, 13095, 13095, 13095, 13095, 13071, 13071, 13071, 13071, 13071, 13071, 13040, 13040, 13040, 13040, 13040, 13040, 13015, 13015, 13015, 13015, 13015, 13015, 13015, 12984, 12984, 12984, 12984, 12984, 12984, 12959, 12959, 12959, 12959, 12959, 12959, 12928, 12928, 12928, 12928, 12928, 12928, 12928, 12904, 12904, 12904, 12904, 12904, 12904, 12873, 12873, 12873, 12873, 12873, 12873, 12848, 12848, 12848, 12848, 12848, 12848, 12848, 12817, 12817, 12817, 12817, 12817, 12817, 12792, 12792, 12792, 12792, 12792, 12792, 12761, 12761, 12761, 12761, 12761, 12761, 12761, 12736, 12736, 12736, 12736, 12736, 12736, 12705, 12705, 12705, 12705, 12705, 12705, 12705, 12681, 12681, 12681, 12681, 12681, 12681, 12650, 12650, 12650, 12650, 12650, 12650, 12625, 12625, 12625, 12625, 12625, 12625, 12625, 12594, 12594, 12594, 12594, 12594, 12594, 12569, 12569, 12569, 12569, 12569, 12569, 12569, 12538, 12538, 12538, 12538, 12538, 12538, 12513, 12513, 12513, 12513, 12513, 12513, 12482, 12482, 12482, 12482, 12482, 12482, 12482, 12457, 12457, 12457, 12457, 12457, 12457, 12426, 12426, 12426, 12426, 12426, 12426, 12426, 12401, 12401, 12401, 12401, 12401, 12401, 12370, 12370, 12370, 12370, 12370, 12370, 12370, 12345, 12345, 12345, 12345, 12345, 12345, 12314, 12314, 12314, 12314, 12314, 12314, 12314, 12289, 12289, 12289, 12289, 12289, 12289, 12258, 12258, 12258, 12258, 12258, 12258, 12258, 12233, 12233, 12233, 12233, 12233, 12233, 12202, 12202, 12202, 12202, 12202, 12202, 12202, 12177, 12177, 12177, 12177, 12177, 12177, 12146, 12146, 12146, 12146, 12146, 12146, 12146, 12121, 12121, 12121, 12121, 12121, 12121, 12090, 12090, 12090, 12090, 12090, 12090, 12090, 12065, 12065, 12065, 12065, 12065, 12065, 12040, 12040, 12040, 12040, 12040, 12040, 12040, 12008, 12008, 12008, 12008, 12008, 12008, 12008, 11983, 11983, 11983, 11983, 11983, 11983, 11952, 11952, 11952, 11952, 11952, 11952, 11952, 11927, 11927, 11927, 11927, 11927, 11927, 11896, 11896, 11896, 11896, 11896, 11896, 11896, 11871, 11871, 11871, 11871, 11871, 11871, 11871, 11840, 11840, 11840, 11840, 11840, 11840, 11815, 11815, 11815, 11815, 11815, 11815, 11815, 11783, 11783, 11783, 11783, 11783, 11783, 11758, 11758, 11758, 11758, 11758, 11758, 11758, 11727, 11727, 11727, 11727, 11727, 11727, 11727, 11702, 11702, 11702, 11702, 11702, 11702, 11670, 11670, 11670, 11670, 11670, 11670, 11670, 11645, 11645, 11645, 11645, 11645, 11645, 11645, 11614, 11614, 11614, 11614, 11614, 11614, 11589, 11589, 11589, 11589, 11589, 11589, 11589, 11558, 11558, 11558, 11558, 11558, 11558, 11558, 11532, 11532, 11532, 11532, 11532, 11532, 11501, 11501, 11501, 11501, 11501, 11501, 11501, 11476, 11476, 11476, 11476, 11476, 11476, 11476, 11444, 11444, 11444, 11444, 11444, 11444, 11444, 11419, 11419, 11419, 11419, 11419, 11419, 11388, 11388, 11388, 11388, 11388, 11388, 11388, 11363, 11363, 11363, 11363, 11363, 11363, 11363, 11331, 11331, 11331, 11331, 11331, 11331, 11331, 11306, 11306, 11306, 11306, 11306, 11306, 11275, 11275, 11275, 11275, 11275, 11275, 11275, 11249, 11249, 11249, 11249, 11249, 11249, 11249, 11218, 11218, 11218, 11218, 11218, 11218, 11218, 11193, 11193, 11193, 11193, 11193, 11193, 11193, 11161, 11161, 11161, 11161, 11161, 11161, 11136, 11136, 11136, 11136, 11136, 11136, 11136, 11104, 11104, 11104, 11104, 11104, 11104, 11104, 11079, 11079, 11079, 11079, 11079, 11079, 11079, 11048, 11048, 11048, 11048, 11048, 11048, 11048, 11022, 11022, 11022, 11022, 11022, 11022, 11022, 10991, 10991, 10991, 10991, 10991, 10991, 10991, 10966, 10966, 10966, 10966, 10966, 10966, 10934, 10934, 10934, 10934, 10934, 10934, 10934, 10909, 10909, 10909, 10909, 10909, 10909, 10909, 10877, 10877, 10877, 10877, 10877, 10877, 10877, 10852, 10852, 10852, 10852, 10852, 10852, 10852, 10820, 10820, 10820, 10820, 10820, 10820, 10820, 10795, 10795, 10795, 10795, 10795, 10795, 10795, 10769, 10769, 10769, 10769, 10769, 10769, 10769, 10738, 10738, 10738, 10738, 10738, 10738, 10738, 10712, 10712, 10712, 10712, 10712, 10712, 10712, 10681, 10681, 10681, 10681, 10681, 10681, 10681, 10655, 10655, 10655, 10655, 10655, 10655, 10655, 10624, 10624, 10624, 10624, 10624, 10624, 10624, 10598, 10598, 10598, 10598, 10598, 10598, 10598, 10567, 10567, 10567, 10567, 10567, 10567, 10567, 10541, 10541, 10541, 10541, 10541, 10541, 10541, 10509, 10509, 10509, 10509, 10509, 10509, 10509, 10484, 10484, 10484, 10484, 10484, 10484, 10484, 10452, 10452, 10452, 10452, 10452, 10452, 10452, 10427, 10427, 10427, 10427, 10427, 10427, 10427, 10395, 10395, 10395, 10395, 10395, 10395, 10395, 10370, 10370, 10370, 10370, 10370, 10370, 10370, 10338, 10338, 10338, 10338, 10338, 10338, 10338, 10312, 10312, 10312, 10312, 10312, 10312, 10312, 10281, 10281, 10281, 10281, 10281, 10281, 10281, 10255, 10255, 10255, 10255, 10255, 10255, 10255, 10255, 10223, 10223, 10223, 10223, 10223, 10223, 10223, 10198, 10198, 10198, 10198, 10198, 10198, 10198, 10166, 10166, 10166, 10166, 10166, 10166, 10166, 10140, 10140, 10140, 10140, 10140, 10140, 10140, 10108, 10108, 10108, 10108, 10108, 10108, 10108, 10083, 10083, 10083, 10083, 10083, 10083, 10083, 10051, 10051, 10051, 10051, 10051, 10051, 10051, 10051, 10025, 10025, 10025, 10025, 10025, 10025, 10025, 9994, 9994, 9994, 9994, 9994, 9994, 9994, 9968, 9968, 9968, 9968, 9968, 9968, 9968, 9936, 9936, 9936, 9936, 9936, 9936, 9936, 9936, 9910, 9910, 9910, 9910, 9910, 9910, 9910, 9878, 9878, 9878, 9878, 9878, 9878, 9878, 9853, 9853, 9853, 9853, 9853, 9853, 9853, 9821, 9821, 9821, 9821, 9821, 9821, 9821, 9821, 9795, 9795, 9795, 9795, 9795, 9795, 9795, 9763, 9763, 9763, 9763, 9763, 9763, 9763, 9738, 9738, 9738, 9738, 9738, 9738, 9738, 9738, 9706, 9706, 9706, 9706, 9706, 9706, 9706, 9680, 9680, 9680, 9680, 9680, 9680, 9680, 9648, 9648, 9648, 9648, 9648, 9648, 9648, 9648, 9622, 9622, 9622, 9622, 9622, 9622, 9622, 9590, 9590, 9590, 9590, 9590, 9590, 9590, 9564, 9564, 9564, 9564, 9564, 9564, 9564, 9564, 9532, 9532, 9532, 9532, 9532, 9532, 9532, 9507, 9507, 9507, 9507, 9507, 9507, 9507, 9481, 9481, 9481, 9481, 9481, 9481, 9481, 9481, 9449, 9449, 9449, 9449, 9449, 9449, 9449, 9423, 9423, 9423, 9423, 9423, 9423, 9423, 9423, 9391, 9391, 9391, 9391, 9391, 9391, 9391, 9365, 9365, 9365, 9365, 9365, 9365, 9365, 9365, 9333, 9333, 9333, 9333, 9333, 9333, 9333, 9307, 9307, 9307, 9307, 9307, 9307, 9307, 9307, 9275, 9275, 9275, 9275, 9275, 9275, 9275, 9249, 9249, 9249, 9249, 9249, 9249, 9249, 9249, 9217, 9217, 9217, 9217, 9217, 9217, 9217, 9191, 9191, 9191, 9191, 9191, 9191, 9191, 9191, 9159, 9159, 9159, 9159, 9159, 9159, 9159, 9133, 9133, 9133, 9133, 9133, 9133, 9133, 9133, 9101, 9101, 9101, 9101, 9101, 9101, 9101, 9075, 9075, 9075, 9075, 9075, 9075, 9075, 9075, 9043, 9043, 9043, 9043, 9043, 9043, 9043, 9017, 9017, 9017, 9017, 9017, 9017, 9017, 9017, 8985, 8985, 8985, 8985, 8985, 8985, 8985, 8985, 8959, 8959, 8959, 8959, 8959, 8959, 8959, 8927, 8927, 8927, 8927, 8927, 8927, 8927, 8927, 8901, 8901, 8901, 8901, 8901, 8901, 8901, 8901, 8868, 8868, 8868, 8868, 8868, 8868, 8868, 8842, 8842, 8842, 8842, 8842, 8842, 8842, 8842, 8810, 8810, 8810, 8810, 8810, 8810, 8810, 8810, 8784, 8784, 8784, 8784, 8784, 8784, 8784, 8752, 8752, 8752, 8752, 8752, 8752, 8752, 8752, 8726, 8726, 8726, 8726, 8726, 8726, 8726, 8726, 8693, 8693, 8693, 8693, 8693, 8693, 8693, 8668, 8668, 8668, 8668, 8668, 8668, 8668, 8668, 8635, 8635, 8635, 8635, 8635, 8635, 8635, 8635, 8609, 8609, 8609, 8609, 8609, 8609, 8609, 8609, 8577, 8577, 8577, 8577, 8577, 8577, 8577, 8577, 8551, 8551, 8551, 8551, 8551, 8551, 8551, 8518, 8518, 8518, 8518, 8518, 8518, 8518, 8518, 8492, 8492, 8492, 8492, 8492, 8492, 8492, 8492, 8460, 8460, 8460, 8460, 8460, 8460, 8460, 8460, 8434, 8434, 8434, 8434, 8434, 8434, 8434, 8434, 8401, 8401, 8401, 8401, 8401, 8401, 8401, 8401, 8375, 8375, 8375, 8375, 8375, 8375, 8375, 8375, 8343, 8343, 8343, 8343, 8343, 8343, 8343, 8316, 8316, 8316, 8316, 8316, 8316, 8316, 8316, 8284, 8284, 8284, 8284, 8284, 8284, 8284, 8284, 8258, 8258, 8258, 8258, 8258, 8258, 8258, 8258, 8232, 8232, 8232, 8232, 8232, 8232, 8232, 8232, 8199, 8199, 8199, 8199, 8199, 8199, 8199, 8199, 8173, 8173, 8173, 8173, 8173, 8173, 8173, 8173, 8140, 8140, 8140, 8140, 8140, 8140, 8140, 8140, 8114, 8114, 8114, 8114, 8114, 8114, 8114, 8114, 8082, 8082, 8082, 8082, 8082, 8082, 8082, 8082, 8056, 8056, 8056, 8056, 8056, 8056, 8056, 8056, 8023, 8023, 8023, 8023, 8023, 8023, 8023, 8023, 7997, 7997, 7997, 7997, 7997, 7997, 7997, 7997, 7964, 7964, 7964, 7964, 7964, 7964, 7964, 7964, 7964, 7938, 7938, 7938, 7938, 7938, 7938, 7938, 7938, 7905, 7905, 7905, 7905, 7905, 7905, 7905, 7905, 7879, 7879, 7879, 7879, 7879, 7879, 7879, 7879, 7846, 7846, 7846, 7846, 7846, 7846, 7846, 7846, 7820, 7820, 7820, 7820, 7820, 7820, 7820, 7820, 7787, 7787, 7787, 7787, 7787, 7787, 7787, 7787, 7761, 7761, 7761, 7761, 7761, 7761, 7761, 7761, 7761, 7728, 7728, 7728, 7728, 7728, 7728, 7728, 7728, 7702, 7702, 7702, 7702, 7702, 7702, 7702, 7702, 7669, 7669, 7669, 7669, 7669, 7669, 7669, 7669, 7643, 7643, 7643, 7643, 7643, 7643, 7643, 7643, 7643, 7610, 7610, 7610, 7610, 7610, 7610, 7610, 7610, 7584, 7584, 7584, 7584, 7584, 7584, 7584, 7584, 7551, 7551, 7551, 7551, 7551, 7551, 7551, 7551, 7551, 7525, 7525, 7525, 7525, 7525, 7525, 7525, 7525, 7492, 7492, 7492, 7492, 7492, 7492, 7492, 7492, 7465, 7465, 7465, 7465, 7465, 7465, 7465, 7465, 7465, 7432, 7432, 7432, 7432, 7432, 7432, 7432, 7432, 7406, 7406, 7406, 7406, 7406, 7406, 7406, 7406, 7373, 7373, 7373, 7373, 7373, 7373, 7373, 7373, 7373, 7347, 7347, 7347, 7347, 7347, 7347, 7347, 7347, 7314, 7314, 7314, 7314, 7314, 7314, 7314, 7314, 7314, 7287, 7287, 7287, 7287, 7287, 7287, 7287, 7287, 7254, 7254, 7254, 7254, 7254, 7254, 7254, 7254, 7254, 7228, 7228, 7228, 7228, 7228, 7228, 7228, 7228, 7195, 7195, 7195, 7195, 7195, 7195, 7195, 7195, 7195, 7169, 7169, 7169, 7169, 7169, 7169, 7169, 7169, 7136, 7136, 7136, 7136, 7136, 7136, 7136, 7136, 7136, 7109, 7109, 7109, 7109, 7109, 7109, 7109, 7109, 7076, 7076, 7076, 7076, 7076, 7076, 7076, 7076, 7076, 7050, 7050, 7050, 7050, 7050, 7050, 7050, 7050, 7050, 7017, 7017, 7017, 7017, 7017, 7017, 7017, 7017, 6990, 6990, 6990, 6990, 6990, 6990, 6990, 6990, 6990, 6957, 6957, 6957, 6957, 6957, 6957, 6957, 6957, 6957, 6931, 6931, 6931, 6931, 6931, 6931, 6931, 6931, 6904, 6904, 6904, 6904, 6904, 6904, 6904, 6904, 6904, 6871, 6871, 6871, 6871, 6871, 6871, 6871, 6871, 6871, 6844, 6844, 6844, 6844, 6844, 6844, 6844, 6844, 6811, 6811, 6811, 6811, 6811, 6811, 6811, 6811, 6811, 6785, 6785, 6785, 6785, 6785, 6785, 6785, 6785, 6785, 6752, 6752, 6752, 6752, 6752, 6752, 6752, 6752, 6752, 6725, 6725, 6725, 6725, 6725, 6725, 6725, 6725, 6725, 6692, 6692, 6692, 6692, 6692, 6692, 6692, 6692, 6692, 6665, 6665, 6665, 6665, 6665, 6665, 6665, 6665, 6632, 6632, 6632, 6632, 6632, 6632, 6632, 6632, 6632, 6605, 6605, 6605, 6605, 6605, 6605, 6605, 6605, 6605, 6572, 6572, 6572, 6572, 6572, 6572, 6572, 6572, 6572, 6545, 6545, 6545, 6545, 6545, 6545, 6545, 6545, 6545, 6512, 6512, 6512, 6512, 6512, 6512, 6512, 6512, 6512, 6486, 6486, 6486, 6486, 6486, 6486, 6486, 6486, 6486, 6452, 6452, 6452, 6452, 6452, 6452, 6452, 6452, 6452, 6426, 6426, 6426, 6426, 6426, 6426, 6426, 6426, 6426, 6392, 6392, 6392, 6392, 6392, 6392, 6392, 6392, 6392, 6366, 6366, 6366, 6366, 6366, 6366, 6366, 6366, 6366, 6332, 6332, 6332, 6332, 6332, 6332, 6332, 6332, 6332, 6305, 6305, 6305, 6305, 6305, 6305, 6305, 6305, 6305, 6272, 6272, 6272, 6272, 6272, 6272, 6272, 6272, 6272, 6272, 6245, 6245, 6245, 6245, 6245, 6245, 6245, 6245, 6245, 6212, 6212, 6212, 6212, 6212, 6212, 6212, 6212, 6212, 6185, 6185, 6185, 6185, 6185, 6185, 6185, 6185, 6185, 6152, 6152, 6152, 6152, 6152, 6152, 6152, 6152, 6152, 6125, 6125, 6125, 6125, 6125, 6125, 6125, 6125, 6125, 6125, 6092, 6092, 6092, 6092, 6092, 6092, 6092, 6092, 6092, 6065, 6065, 6065, 6065, 6065, 6065, 6065, 6065, 6065, 6031, 6031, 6031, 6031, 6031, 6031, 6031, 6031, 6031, 6005, 6005, 6005, 6005, 6005, 6005, 6005, 6005, 6005, 6005, 5971, 5971, 5971, 5971, 5971, 5971, 5971, 5971, 5971, 5944, 5944, 5944, 5944, 5944, 5944, 5944, 5944, 5944, 5944, 5911, 5911, 5911, 5911, 5911, 5911, 5911, 5911, 5911, 5884, 5884, 5884, 5884, 5884, 5884, 5884, 5884, 5884, 5850, 5850, 5850, 5850, 5850, 5850, 5850, 5850, 5850, 5850, 5823, 5823, 5823, 5823, 5823, 5823, 5823, 5823, 5823, 5790, 5790, 5790, 5790, 5790, 5790, 5790, 5790, 5790, 5790, 5763, 5763, 5763, 5763, 5763, 5763, 5763, 5763, 5763, 5729, 5729, 5729, 5729, 5729, 5729, 5729, 5729, 5729, 5729, 5702, 5702, 5702, 5702, 5702, 5702, 5702, 5702, 5702, 5702, 5669, 5669, 5669, 5669, 5669, 5669, 5669, 5669, 5669, 5642, 5642, 5642, 5642, 5642, 5642, 5642, 5642, 5642, 5642, 5608, 5608, 5608, 5608, 5608, 5608, 5608, 5608, 5608, 5608, 5581, 5581, 5581, 5581, 5581, 5581, 5581, 5581, 5581, 5554, 5554, 5554, 5554, 5554, 5554, 5554, 5554, 5554, 5554, 5521, 5521, 5521, 5521, 5521, 5521, 5521, 5521, 5521, 5521, 5494, 5494, 5494, 5494, 5494, 5494, 5494, 5494, 5494, 5494, 5460, 5460, 5460, 5460, 5460, 5460, 5460, 5460, 5460, 5433, 5433, 5433, 5433, 5433, 5433, 5433, 5433, 5433, 5433, 5399, 5399, 5399, 5399, 5399, 5399, 5399, 5399, 5399, 5399, 5372, 5372, 5372, 5372, 5372, 5372, 5372, 5372, 5372, 5372, 5338, 5338, 5338, 5338, 5338, 5338, 5338, 5338, 5338, 5338, 5311, 5311, 5311, 5311, 5311, 5311, 5311, 5311, 5311, 5311, 5278, 5278, 5278, 5278, 5278, 5278, 5278, 5278, 5278, 5278, 5250, 5250, 5250, 5250, 5250, 5250, 5250, 5250, 5250, 5250, 5217, 5217, 5217, 5217, 5217, 5217, 5217, 5217, 5217, 5217, 5190, 5190, 5190, 5190, 5190, 5190, 5190, 5190, 5190, 5190, 5156, 5156, 5156, 5156, 5156, 5156, 5156, 5156, 5156, 5156, 5129, 5129, 5129, 5129, 5129, 5129, 5129, 5129, 5129, 5129, 5095, 5095, 5095, 5095, 5095, 5095, 5095, 5095, 5095, 5095, 5068, 5068, 5068, 5068, 5068, 5068, 5068, 5068, 5068, 5068, 5034, 5034, 5034, 5034, 5034, 5034, 5034, 5034, 5034, 5034, 5034, 5007, 5007, 5007, 5007, 5007, 5007, 5007, 5007, 5007, 5007, 4973, 4973, 4973, 4973, 4973, 4973, 4973, 4973, 4973, 4973, 4945, 4945, 4945, 4945, 4945, 4945, 4945, 4945, 4945, 4945, 4945, 4912, 4912, 4912, 4912, 4912, 4912, 4912, 4912, 4912, 4912, 4884, 4884, 4884, 4884, 4884, 4884, 4884, 4884, 4884, 4884, 4850, 4850, 4850, 4850, 4850, 4850, 4850, 4850, 4850, 4850, 4850, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4789, 4789, 4789, 4789, 4789, 4789, 4789, 4789, 4789, 4789, 4789, 4762, 4762, 4762, 4762, 4762, 4762, 4762, 4762, 4762, 4762, 4728, 4728, 4728, 4728, 4728, 4728, 4728, 4728, 4728, 4728, 4728, 4701, 4701, 4701, 4701, 4701, 4701, 4701, 4701, 4701, 4701, 4667, 4667, 4667, 4667, 4667, 4667, 4667, 4667, 4667, 4667, 4667, 4639, 4639, 4639, 4639, 4639, 4639, 4639, 4639, 4639, 4639, 4605, 4605, 4605, 4605, 4605, 4605, 4605, 4605, 4605, 4605, 4605, 4578, 4578, 4578, 4578, 4578, 4578, 4578, 4578, 4578, 4578, 4578, 4544, 4544, 4544, 4544, 4544, 4544, 4544, 4544, 4544, 4544, 4544, 4516, 4516, 4516, 4516, 4516, 4516, 4516, 4516, 4516, 4516, 4482, 4482, 4482, 4482, 4482, 4482, 4482, 4482, 4482, 4482, 4482, 4455, 4455, 4455, 4455, 4455, 4455, 4455, 4455, 4455, 4455, 4455, 4421, 4421, 4421, 4421, 4421, 4421, 4421, 4421, 4421, 4421, 4421, 4393, 4393, 4393, 4393, 4393, 4393, 4393, 4393, 4393, 4393, 4393, 4359, 4359, 4359, 4359, 4359, 4359, 4359, 4359, 4359, 4359, 4359, 4332, 4332, 4332, 4332, 4332, 4332, 4332, 4332, 4332, 4332, 4332, 4298, 4298, 4298, 4298, 4298, 4298, 4298, 4298, 4298, 4298, 4298, 4270, 4270, 4270, 4270, 4270, 4270, 4270, 4270, 4270, 4270, 4270, 4236, 4236, 4236, 4236, 4236, 4236, 4236, 4236, 4236, 4236, 4236, 4209, 4209, 4209, 4209, 4209, 4209, 4209, 4209, 4209, 4209, 4209, 4209, 4181, 4181, 4181, 4181, 4181, 4181, 4181, 4181, 4181, 4181, 4181, 4147, 4147, 4147, 4147, 4147, 4147, 4147, 4147, 4147, 4147, 4147, 4119, 4119, 4119, 4119, 4119, 4119, 4119, 4119, 4119, 4119, 4119, 4085, 4085, 4085, 4085, 4085, 4085, 4085, 4085, 4085, 4085, 4085, 4085, 4058, 4058, 4058, 4058, 4058, 4058, 4058, 4058, 4058, 4058, 4058, 4023, 4023, 4023, 4023, 4023, 4023, 4023, 4023, 4023, 4023, 4023, 4023, 3996, 3996, 3996, 3996, 3996, 3996, 3996, 3996, 3996, 3996, 3996, 3961, 3961, 3961, 3961, 3961, 3961, 3961, 3961, 3961, 3961, 3961, 3961, 3934, 3934, 3934, 3934, 3934, 3934, 3934, 3934, 3934, 3934, 3934, 3899, 3899, 3899, 3899, 3899, 3899, 3899, 3899, 3899, 3899, 3899, 3899, 3872, 3872, 3872, 3872, 3872, 3872, 3872, 3872, 3872, 3872, 3872, 3837, 3837, 3837, 3837, 3837, 3837, 3837, 3837, 3837, 3837, 3837, 3837, 3810, 3810, 3810, 3810, 3810, 3810, 3810, 3810, 3810, 3810, 3810, 3810, 3775, 3775, 3775, 3775, 3775, 3775, 3775, 3775, 3775, 3775, 3775, 3775, 3748, 3748, 3748, 3748, 3748, 3748, 3748, 3748, 3748, 3748, 3748, 3748, 3713, 3713, 3713, 3713, 3713, 3713, 3713, 3713, 3713, 3713, 3713, 3713, 3686, 3686, 3686, 3686, 3686, 3686, 3686, 3686, 3686, 3686, 3686, 3686, 3651, 3651, 3651, 3651, 3651, 3651, 3651, 3651, 3651, 3651, 3651, 3651, 3624, 3624, 3624, 3624, 3624, 3624, 3624, 3624, 3624, 3624, 3624, 3624, 3589, 3589, 3589, 3589, 3589, 3589, 3589, 3589, 3589, 3589, 3589, 3589, 3561, 3561, 3561, 3561, 3561, 3561, 3561, 3561, 3561, 3561, 3561, 3561, 3527, 3527, 3527, 3527, 3527, 3527, 3527, 3527, 3527, 3527, 3527, 3527, 3499, 3499, 3499, 3499, 3499, 3499, 3499, 3499, 3499, 3499, 3499, 3499, 3465, 3465, 3465, 3465, 3465, 3465, 3465, 3465, 3465, 3465, 3465, 3465, 3465, 3437, 3437, 3437, 3437, 3437, 3437, 3437, 3437, 3437, 3437, 3437, 3437, 3402, 3402, 3402, 3402, 3402, 3402, 3402, 3402, 3402, 3402, 3402, 3402, 3402, 3374, 3374, 3374, 3374, 3374, 3374, 3374, 3374, 3374, 3374, 3374, 3374, 3340, 3340, 3340, 3340, 3340, 3340, 3340, 3340, 3340, 3340, 3340, 3340, 3340, 3312, 3312, 3312, 3312, 3312, 3312, 3312, 3312, 3312, 3312, 3312, 3312, 3277, 3277, 3277, 3277, 3277, 3277, 3277, 3277, 3277, 3277, 3277, 3277, 3277, 3250, 3250, 3250, 3250, 3250, 3250, 3250, 3250, 3250, 3250, 3250, 3250, 3250, 3215, 3215, 3215, 3215, 3215, 3215, 3215, 3215, 3215, 3215, 3215, 3215, 3215, 3187, 3187, 3187, 3187, 3187, 3187, 3187, 3187, 3187, 3187, 3187, 3187, 3152, 3152, 3152, 3152, 3152, 3152, 3152, 3152, 3152, 3152, 3152, 3152, 3152, 3125, 3125, 3125, 3125, 3125, 3125, 3125, 3125, 3125, 3125, 3125, 3125, 3125, 3090, 3090, 3090, 3090, 3090, 3090, 3090, 3090, 3090, 3090, 3090, 3090, 3090, 3062, 3062, 3062, 3062, 3062, 3062, 3062, 3062, 3062, 3062, 3062, 3062, 3062, 3062, 3027, 3027, 3027, 3027, 3027, 3027, 3027, 3027, 3027, 3027, 3027, 3027, 3027, 2999, 2999, 2999, 2999, 2999, 2999, 2999, 2999, 2999, 2999, 2999, 2999, 2999, 2964, 2964, 2964, 2964, 2964, 2964, 2964, 2964, 2964, 2964, 2964, 2964, 2964, 2937, 2937, 2937, 2937, 2937, 2937, 2937, 2937, 2937, 2937, 2937, 2937, 2937, 2937, 2902, 2902, 2902, 2902, 2902, 2902, 2902, 2902, 2902, 2902, 2902, 2902, 2902, 2874, 2874, 2874, 2874, 2874, 2874, 2874, 2874, 2874, 2874, 2874, 2874, 2874, 2874, 2846, 2846, 2846, 2846, 2846, 2846, 2846, 2846, 2846, 2846, 2846, 2846, 2846, 2846, 2811, 2811, 2811, 2811, 2811, 2811, 2811, 2811, 2811, 2811, 2811, 2811, 2811, 2783, 2783, 2783, 2783, 2783, 2783, 2783, 2783, 2783, 2783, 2783, 2783, 2783, 2783, 2748, 2748, 2748, 2748, 2748, 2748, 2748, 2748, 2748, 2748, 2748, 2748, 2748, 2748, 2720, 2720, 2720, 2720, 2720, 2720, 2720, 2720, 2720, 2720, 2720, 2720, 2720, 2720, 2685, 2685, 2685, 2685, 2685, 2685, 2685, 2685, 2685, 2685, 2685, 2685, 2685, 2685, 2657, 2657, 2657, 2657, 2657, 2657, 2657, 2657, 2657, 2657, 2657, 2657, 2657, 2657, 2622, 2622, 2622, 2622, 2622, 2622, 2622, 2622, 2622, 2622, 2622, 2622, 2622, 2622, 2594, 2594, 2594, 2594, 2594, 2594, 2594, 2594, 2594, 2594, 2594, 2594, 2594, 2594, 2594, 2559, 2559, 2559, 2559, 2559, 2559, 2559, 2559, 2559, 2559, 2559, 2559, 2559, 2559, 2531, 2531, 2531, 2531, 2531, 2531, 2531, 2531, 2531, 2531, 2531, 2531, 2531, 2531, 2496, 2496, 2496, 2496, 2496, 2496, 2496, 2496, 2496, 2496, 2496, 2496, 2496, 2496, 2496, 2468, 2468, 2468, 2468, 2468, 2468, 2468, 2468, 2468, 2468, 2468, 2468, 2468, 2468, 2468, 2433, 2433, 2433, 2433, 2433, 2433, 2433, 2433, 2433, 2433, 2433, 2433, 2433, 2433, 2405, 2405, 2405, 2405, 2405, 2405, 2405, 2405, 2405, 2405, 2405, 2405, 2405, 2405, 2405, 2370, 2370, 2370, 2370, 2370, 2370, 2370, 2370, 2370, 2370, 2370, 2370, 2370, 2370, 2370, 2342, 2342, 2342, 2342, 2342, 2342, 2342, 2342, 2342, 2342, 2342, 2342, 2342, 2342, 2342, 2307, 2307, 2307, 2307, 2307, 2307, 2307, 2307, 2307, 2307, 2307, 2307, 2307, 2307, 2307, 2278, 2278, 2278, 2278, 2278, 2278, 2278, 2278, 2278, 2278, 2278, 2278, 2278, 2278, 2278, 2278, 2243, 2243, 2243, 2243, 2243, 2243, 2243, 2243, 2243, 2243, 2243, 2243, 2243, 2243, 2243, 2215, 2215, 2215, 2215, 2215, 2215, 2215, 2215, 2215, 2215, 2215, 2215, 2215, 2215, 2215, 2180, 2180, 2180, 2180, 2180, 2180, 2180, 2180, 2180, 2180, 2180, 2180, 2180, 2180, 2180, 2180, 2152, 2152, 2152, 2152, 2152, 2152, 2152, 2152, 2152, 2152, 2152, 2152, 2152, 2152, 2152, 2152, 2116, 2116, 2116, 2116, 2116, 2116, 2116, 2116, 2116, 2116, 2116, 2116, 2116, 2116, 2116, 2088, 2088, 2088, 2088, 2088, 2088, 2088, 2088, 2088, 2088, 2088, 2088, 2088, 2088, 2088, 2088, 2053, 2053, 2053, 2053, 2053, 2053, 2053, 2053, 2053, 2053, 2053, 2053, 2053, 2053, 2053, 2053, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 1989, 1989, 1989, 1989, 1989, 1989, 1989, 1989, 1989, 1989, 1989, 1989, 1989, 1989, 1989, 1989, 1961, 1961, 1961, 1961, 1961, 1961, 1961, 1961, 1961, 1961, 1961, 1961, 1961, 1961, 1961, 1961, 1926, 1926, 1926, 1926, 1926, 1926, 1926, 1926, 1926, 1926, 1926, 1926, 1926, 1926, 1926, 1926, 1926, 1898, 1898, 1898, 1898, 1898, 1898, 1898, 1898, 1898, 1898, 1898, 1898, 1898, 1898, 1898, 1898, 1898, 1862, 1862, 1862, 1862, 1862, 1862, 1862, 1862, 1862, 1862, 1862, 1862, 1862, 1862, 1862, 1862, 1862, 1834, 1834, 1834, 1834, 1834, 1834, 1834, 1834, 1834, 1834, 1834, 1834, 1834, 1834, 1834, 1834, 1834, 1799, 1799, 1799, 1799, 1799, 1799, 1799, 1799, 1799, 1799, 1799, 1799, 1799, 1799, 1799, 1799, 1799, 1770, 1770, 1770, 1770, 1770, 1770, 1770, 1770, 1770, 1770, 1770, 1770, 1770, 1770, 1770, 1770, 1770, 1735, 1735, 1735, 1735, 1735, 1735, 1735, 1735, 1735, 1735, 1735, 1735, 1735, 1735, 1735, 1735, 1735, 1735, 1707, 1707, 1707, 1707, 1707, 1707, 1707, 1707, 1707, 1707, 1707, 1707, 1707, 1707, 1707, 1707, 1707, 1671, 1671, 1671, 1671, 1671, 1671, 1671, 1671, 1671, 1671, 1671, 1671, 1671, 1671, 1671, 1671, 1671, 1671, 1643, 1643, 1643, 1643, 1643, 1643, 1643, 1643, 1643, 1643, 1643, 1643, 1643, 1643, 1643, 1643, 1643, 1643, 1607, 1607, 1607, 1607, 1607, 1607, 1607, 1607, 1607, 1607, 1607, 1607, 1607, 1607, 1607, 1607, 1607, 1607, 1579, 1579, 1579, 1579, 1579, 1579, 1579, 1579, 1579, 1579, 1579, 1579, 1579, 1579, 1579, 1579, 1579, 1579, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70421, 70421, 70421, 70421, 70421, 70421, 70421, 70421, 70421, 70421, 70421, 70421, 70421, 70421, 70421, 70421, 70421, 70421, 70393, 70393, 70393, 70393, 70393, 70393, 70393, 70393, 70393, 70393, 70393, 70393, 70393, 70393, 70393, 70393, 70393, 70393, 70357, 70357, 70357, 70357, 70357, 70357, 70357, 70357, 70357, 70357, 70357, 70357, 70357, 70357, 70357, 70357, 70357, 70357, 70329, 70329, 70329, 70329, 70329, 70329, 70329, 70329, 70329, 70329, 70329, 70329, 70329, 70329, 70329, 70329, 70329, 70329, 70293, 70293, 70293, 70293, 70293, 70293, 70293, 70293, 70293, 70293, 70293, 70293, 70293, 70293, 70293, 70293, 70293, 70265, 70265, 70265, 70265, 70265, 70265, 70265, 70265, 70265, 70265, 70265, 70265, 70265, 70265, 70265, 70265, 70265, 70265, 70230, 70230, 70230, 70230, 70230, 70230, 70230, 70230, 70230, 70230, 70230, 70230, 70230, 70230, 70230, 70230, 70230, 70201, 70201, 70201, 70201, 70201, 70201, 70201, 70201, 70201, 70201, 70201, 70201, 70201, 70201, 70201, 70201, 70201, 70166, 70166, 70166, 70166, 70166, 70166, 70166, 70166, 70166, 70166, 70166, 70166, 70166, 70166, 70166, 70166, 70166, 70138, 70138, 70138, 70138, 70138, 70138, 70138, 70138, 70138, 70138, 70138, 70138, 70138, 70138, 70138, 70138, 70138, 70102, 70102, 70102, 70102, 70102, 70102, 70102, 70102, 70102, 70102, 70102, 70102, 70102, 70102, 70102, 70102, 70102, 70074, 70074, 70074, 70074, 70074, 70074, 70074, 70074, 70074, 70074, 70074, 70074, 70074, 70074, 70074, 70074, 70074, 70039, 70039, 70039, 70039, 70039, 70039, 70039, 70039, 70039, 70039, 70039, 70039, 70039, 70039, 70039, 70039, 70011, 70011, 70011, 70011, 70011, 70011, 70011, 70011, 70011, 70011, 70011, 70011, 70011, 70011, 70011, 70011, 69975, 69975, 69975, 69975, 69975, 69975, 69975, 69975, 69975, 69975, 69975, 69975, 69975, 69975, 69975, 69975, 69975, 69947, 69947, 69947, 69947, 69947, 69947, 69947, 69947, 69947, 69947, 69947, 69947, 69947, 69947, 69947, 69947, 69912, 69912, 69912, 69912, 69912, 69912, 69912, 69912, 69912, 69912, 69912, 69912, 69912, 69912, 69912, 69912, 69884, 69884, 69884, 69884, 69884, 69884, 69884, 69884, 69884, 69884, 69884, 69884, 69884, 69884, 69884, 69848, 69848, 69848, 69848, 69848, 69848, 69848, 69848, 69848, 69848, 69848, 69848, 69848, 69848, 69848, 69848, 69820, 69820, 69820, 69820, 69820, 69820, 69820, 69820, 69820, 69820, 69820, 69820, 69820, 69820, 69820, 69820, 69785, 69785, 69785, 69785, 69785, 69785, 69785, 69785, 69785, 69785, 69785, 69785, 69785, 69785, 69785, 69757, 69757, 69757, 69757, 69757, 69757, 69757, 69757, 69757, 69757, 69757, 69757, 69757, 69757, 69757, 69722, 69722, 69722, 69722, 69722, 69722, 69722, 69722, 69722, 69722, 69722, 69722, 69722, 69722, 69722, 69722, 69693, 69693, 69693, 69693, 69693, 69693, 69693, 69693, 69693, 69693, 69693, 69693, 69693, 69693, 69693, 69658, 69658, 69658, 69658, 69658, 69658, 69658, 69658, 69658, 69658, 69658, 69658, 69658, 69658, 69658, 69630, 69630, 69630, 69630, 69630, 69630, 69630, 69630, 69630, 69630, 69630, 69630, 69630, 69630, 69630, 69595, 69595, 69595, 69595, 69595, 69595, 69595, 69595, 69595, 69595, 69595, 69595, 69595, 69595, 69595, 69567, 69567, 69567, 69567, 69567, 69567, 69567, 69567, 69567, 69567, 69567, 69567, 69567, 69567, 69532, 69532, 69532, 69532, 69532, 69532, 69532, 69532, 69532, 69532, 69532, 69532, 69532, 69532, 69532, 69504, 69504, 69504, 69504, 69504, 69504, 69504, 69504, 69504, 69504, 69504, 69504, 69504, 69504, 69504, 69469, 69469, 69469, 69469, 69469, 69469, 69469, 69469, 69469, 69469, 69469, 69469, 69469, 69469, 69441, 69441, 69441, 69441, 69441, 69441, 69441, 69441, 69441, 69441, 69441, 69441, 69441, 69441, 69406, 69406, 69406, 69406, 69406, 69406, 69406, 69406, 69406, 69406, 69406, 69406, 69406, 69406, 69406, 69378, 69378, 69378, 69378, 69378, 69378, 69378, 69378, 69378, 69378, 69378, 69378, 69378, 69378, 69343, 69343, 69343, 69343, 69343, 69343, 69343, 69343, 69343, 69343, 69343, 69343, 69343, 69343, 69315, 69315, 69315, 69315, 69315, 69315, 69315, 69315, 69315, 69315, 69315, 69315, 69315, 69315, 69280, 69280, 69280, 69280, 69280, 69280, 69280, 69280, 69280, 69280, 69280, 69280, 69280, 69280, 69252, 69252, 69252, 69252, 69252, 69252, 69252, 69252, 69252, 69252, 69252, 69252, 69252, 69252, 69217, 69217, 69217, 69217, 69217, 69217, 69217, 69217, 69217, 69217, 69217, 69217, 69217, 69217, 69189, 69189, 69189, 69189, 69189, 69189, 69189, 69189, 69189, 69189, 69189, 69189, 69189, 69154, 69154, 69154, 69154, 69154, 69154, 69154, 69154, 69154, 69154, 69154, 69154, 69154, 69154, 69126, 69126, 69126, 69126, 69126, 69126, 69126, 69126, 69126, 69126, 69126, 69126, 69126, 69126, 69098, 69098, 69098, 69098, 69098, 69098, 69098, 69098, 69098, 69098, 69098, 69098, 69098, 69063, 69063, 69063, 69063, 69063, 69063, 69063, 69063, 69063, 69063, 69063, 69063, 69063, 69063, 69036, 69036, 69036, 69036, 69036, 69036, 69036, 69036, 69036, 69036, 69036, 69036, 69036, 69001, 69001, 69001, 69001, 69001, 69001, 69001, 69001, 69001, 69001, 69001, 69001, 69001, 68973, 68973, 68973, 68973, 68973, 68973, 68973, 68973, 68973, 68973, 68973, 68973, 68973, 68938, 68938, 68938, 68938, 68938, 68938, 68938, 68938, 68938, 68938, 68938, 68938, 68938, 68938, 68910, 68910, 68910, 68910, 68910, 68910, 68910, 68910, 68910, 68910, 68910, 68910, 68910, 68875, 68875, 68875, 68875, 68875, 68875, 68875, 68875, 68875, 68875, 68875, 68875, 68875, 68848, 68848, 68848, 68848, 68848, 68848, 68848, 68848, 68848, 68848, 68848, 68848, 68848, 68813, 68813, 68813, 68813, 68813, 68813, 68813, 68813, 68813, 68813, 68813, 68813, 68785, 68785, 68785, 68785, 68785, 68785, 68785, 68785, 68785, 68785, 68785, 68785, 68785, 68750, 68750, 68750, 68750, 68750, 68750, 68750, 68750, 68750, 68750, 68750, 68750, 68750, 68723, 68723, 68723, 68723, 68723, 68723, 68723, 68723, 68723, 68723, 68723, 68723, 68723, 68688, 68688, 68688, 68688, 68688, 68688, 68688, 68688, 68688, 68688, 68688, 68688, 68660, 68660, 68660, 68660, 68660, 68660, 68660, 68660, 68660, 68660, 68660, 68660, 68660, 68626, 68626, 68626, 68626, 68626, 68626, 68626, 68626, 68626, 68626, 68626, 68626, 68598, 68598, 68598, 68598, 68598, 68598, 68598, 68598, 68598, 68598, 68598, 68598, 68598, 68563, 68563, 68563, 68563, 68563, 68563, 68563, 68563, 68563, 68563, 68563, 68563, 68535, 68535, 68535, 68535, 68535, 68535, 68535, 68535, 68535, 68535, 68535, 68535, 68535, 68501, 68501, 68501, 68501, 68501, 68501, 68501, 68501, 68501, 68501, 68501, 68501, 68473, 68473, 68473, 68473, 68473, 68473, 68473, 68473, 68473, 68473, 68473, 68473, 68439, 68439, 68439, 68439, 68439, 68439, 68439, 68439, 68439, 68439, 68439, 68439, 68411, 68411, 68411, 68411, 68411, 68411, 68411, 68411, 68411, 68411, 68411, 68411, 68376, 68376, 68376, 68376, 68376, 68376, 68376, 68376, 68376, 68376, 68376, 68376, 68349, 68349, 68349, 68349, 68349, 68349, 68349, 68349, 68349, 68349, 68349, 68349, 68314, 68314, 68314, 68314, 68314, 68314, 68314, 68314, 68314, 68314, 68314, 68314, 68287, 68287, 68287, 68287, 68287, 68287, 68287, 68287, 68287, 68287, 68287, 68287, 68252, 68252, 68252, 68252, 68252, 68252, 68252, 68252, 68252, 68252, 68252, 68252, 68225, 68225, 68225, 68225, 68225, 68225, 68225, 68225, 68225, 68225, 68225, 68225, 68190, 68190, 68190, 68190, 68190, 68190, 68190, 68190, 68190, 68190, 68190, 68190, 68163, 68163, 68163, 68163, 68163, 68163, 68163, 68163, 68163, 68163, 68163, 68163, 68128, 68128, 68128, 68128, 68128, 68128, 68128, 68128, 68128, 68128, 68128, 68101, 68101, 68101, 68101, 68101, 68101, 68101, 68101, 68101, 68101, 68101, 68101, 68066, 68066, 68066, 68066, 68066, 68066, 68066, 68066, 68066, 68066, 68066, 68039, 68039, 68039, 68039, 68039, 68039, 68039, 68039, 68039, 68039, 68039, 68039, 68004, 68004, 68004, 68004, 68004, 68004, 68004, 68004, 68004, 68004, 68004, 67977, 67977, 67977, 67977, 67977, 67977, 67977, 67977, 67977, 67977, 67977, 67977, 67942, 67942, 67942, 67942, 67942, 67942, 67942, 67942, 67942, 67942, 67942, 67915, 67915, 67915, 67915, 67915, 67915, 67915, 67915, 67915, 67915, 67915, 67915, 67881, 67881, 67881, 67881, 67881, 67881, 67881, 67881, 67881, 67881, 67881, 67853, 67853, 67853, 67853, 67853, 67853, 67853, 67853, 67853, 67853, 67853, 67819, 67819, 67819, 67819, 67819, 67819, 67819, 67819, 67819, 67819, 67819, 67791, 67791, 67791, 67791, 67791, 67791, 67791, 67791, 67791, 67791, 67791, 67791, 67764, 67764, 67764, 67764, 67764, 67764, 67764, 67764, 67764, 67764, 67764, 67730, 67730, 67730, 67730, 67730, 67730, 67730, 67730, 67730, 67730, 67730, 67702, 67702, 67702, 67702, 67702, 67702, 67702, 67702, 67702, 67702, 67702, 67668, 67668, 67668, 67668, 67668, 67668, 67668, 67668, 67668, 67668, 67668, 67641, 67641, 67641, 67641, 67641, 67641, 67641, 67641, 67641, 67641, 67641, 67607, 67607, 67607, 67607, 67607, 67607, 67607, 67607, 67607, 67607, 67607, 67579, 67579, 67579, 67579, 67579, 67579, 67579, 67579, 67579, 67579, 67579, 67545, 67545, 67545, 67545, 67545, 67545, 67545, 67545, 67545, 67545, 67545, 67518, 67518, 67518, 67518, 67518, 67518, 67518, 67518, 67518, 67518, 67518, 67484, 67484, 67484, 67484, 67484, 67484, 67484, 67484, 67484, 67484, 67456, 67456, 67456, 67456, 67456, 67456, 67456, 67456, 67456, 67456, 67456, 67422, 67422, 67422, 67422, 67422, 67422, 67422, 67422, 67422, 67422, 67422, 67395, 67395, 67395, 67395, 67395, 67395, 67395, 67395, 67395, 67395, 67395, 67361, 67361, 67361, 67361, 67361, 67361, 67361, 67361, 67361, 67361, 67333, 67333, 67333, 67333, 67333, 67333, 67333, 67333, 67333, 67333, 67333, 67299, 67299, 67299, 67299, 67299, 67299, 67299, 67299, 67299, 67299, 67272, 67272, 67272, 67272, 67272, 67272, 67272, 67272, 67272, 67272, 67272, 67238, 67238, 67238, 67238, 67238, 67238, 67238, 67238, 67238, 67238, 67211, 67211, 67211, 67211, 67211, 67211, 67211, 67211, 67211, 67211, 67211, 67177, 67177, 67177, 67177, 67177, 67177, 67177, 67177, 67177, 67177, 67150, 67150, 67150, 67150, 67150, 67150, 67150, 67150, 67150, 67150, 67150, 67116, 67116, 67116, 67116, 67116, 67116, 67116, 67116, 67116, 67116, 67088, 67088, 67088, 67088, 67088, 67088, 67088, 67088, 67088, 67088, 67055, 67055, 67055, 67055, 67055, 67055, 67055, 67055, 67055, 67055, 67055, 67027, 67027, 67027, 67027, 67027, 67027, 67027, 67027, 67027, 67027, 66993, 66993, 66993, 66993, 66993, 66993, 66993, 66993, 66993, 66993, 66966, 66966, 66966, 66966, 66966, 66966, 66966, 66966, 66966, 66966, 66966, 66932, 66932, 66932, 66932, 66932, 66932, 66932, 66932, 66932, 66932, 66905, 66905, 66905, 66905, 66905, 66905, 66905, 66905, 66905, 66905, 66871, 66871, 66871, 66871, 66871, 66871, 66871, 66871, 66871, 66871, 66844, 66844, 66844, 66844, 66844, 66844, 66844, 66844, 66844, 66844, 66810, 66810, 66810, 66810, 66810, 66810, 66810, 66810, 66810, 66810, 66783, 66783, 66783, 66783, 66783, 66783, 66783, 66783, 66783, 66783, 66750, 66750, 66750, 66750, 66750, 66750, 66750, 66750, 66750, 66750, 66722, 66722, 66722, 66722, 66722, 66722, 66722, 66722, 66722, 66722, 66689, 66689, 66689, 66689, 66689, 66689, 66689, 66689, 66689, 66689, 66662, 66662, 66662, 66662, 66662, 66662, 66662, 66662, 66662, 66662, 66628, 66628, 66628, 66628, 66628, 66628, 66628, 66628, 66628, 66628, 66601, 66601, 66601, 66601, 66601, 66601, 66601, 66601, 66601, 66601, 66567, 66567, 66567, 66567, 66567, 66567, 66567, 66567, 66567, 66567, 66540, 66540, 66540, 66540, 66540, 66540, 66540, 66540, 66540, 66506, 66506, 66506, 66506, 66506, 66506, 66506, 66506, 66506, 66506, 66479, 66479, 66479, 66479, 66479, 66479, 66479, 66479, 66479, 66479, 66446, 66446, 66446, 66446, 66446, 66446, 66446, 66446, 66446, 66446, 66419, 66419, 66419, 66419, 66419, 66419, 66419, 66419, 66419, 66392, 66392, 66392, 66392, 66392, 66392, 66392, 66392, 66392, 66392, 66358, 66358, 66358, 66358, 66358, 66358, 66358, 66358, 66358, 66358, 66331, 66331, 66331, 66331, 66331, 66331, 66331, 66331, 66331, 66298, 66298, 66298, 66298, 66298, 66298, 66298, 66298, 66298, 66298, 66271, 66271, 66271, 66271, 66271, 66271, 66271, 66271, 66271, 66271, 66237, 66237, 66237, 66237, 66237, 66237, 66237, 66237, 66237, 66210, 66210, 66210, 66210, 66210, 66210, 66210, 66210, 66210, 66210, 66177, 66177, 66177, 66177, 66177, 66177, 66177, 66177, 66177, 66150, 66150, 66150, 66150, 66150, 66150, 66150, 66150, 66150, 66150, 66116, 66116, 66116, 66116, 66116, 66116, 66116, 66116, 66116, 66089, 66089, 66089, 66089, 66089, 66089, 66089, 66089, 66089, 66056, 66056, 66056, 66056, 66056, 66056, 66056, 66056, 66056, 66056, 66029, 66029, 66029, 66029, 66029, 66029, 66029, 66029, 66029, 65995, 65995, 65995, 65995, 65995, 65995, 65995, 65995, 65995, 65995, 65969, 65969, 65969, 65969, 65969, 65969, 65969, 65969, 65969, 65935, 65935, 65935, 65935, 65935, 65935, 65935, 65935, 65935, 65908, 65908, 65908, 65908, 65908, 65908, 65908, 65908, 65908, 65875, 65875, 65875, 65875, 65875, 65875, 65875, 65875, 65875, 65875, 65848, 65848, 65848, 65848, 65848, 65848, 65848, 65848, 65848, 65815, 65815, 65815, 65815, 65815, 65815, 65815, 65815, 65815, 65788, 65788, 65788, 65788, 65788, 65788, 65788, 65788, 65788, 65755, 65755, 65755, 65755, 65755, 65755, 65755, 65755, 65755, 65728, 65728, 65728, 65728, 65728, 65728, 65728, 65728, 65728, 65728, 65695, 65695, 65695, 65695, 65695, 65695, 65695, 65695, 65695, 65668, 65668, 65668, 65668, 65668, 65668, 65668, 65668, 65668, 65634, 65634, 65634, 65634, 65634, 65634, 65634, 65634, 65634, 65608, 65608, 65608, 65608, 65608, 65608, 65608, 65608, 65608, 65574, 65574, 65574, 65574, 65574, 65574, 65574, 65574, 65574, 65548, 65548, 65548, 65548, 65548, 65548, 65548, 65548, 65548, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65455, 65455, 65455, 65455, 65455, 65455, 65455, 65455, 65455, 65428, 65428, 65428, 65428, 65428, 65428, 65428, 65428, 65428, 65395, 65395, 65395, 65395, 65395, 65395, 65395, 65395, 65395, 65368, 65368, 65368, 65368, 65368, 65368, 65368, 65368, 65368, 65335, 65335, 65335, 65335, 65335, 65335, 65335, 65335, 65308, 65308, 65308, 65308, 65308, 65308, 65308, 65308, 65308, 65275, 65275, 65275, 65275, 65275, 65275, 65275, 65275, 65275, 65248, 65248, 65248, 65248, 65248, 65248, 65248, 65248, 65248, 65215, 65215, 65215, 65215, 65215, 65215, 65215, 65215, 65215, 65189, 65189, 65189, 65189, 65189, 65189, 65189, 65189, 65189, 65156, 65156, 65156, 65156, 65156, 65156, 65156, 65156, 65129, 65129, 65129, 65129, 65129, 65129, 65129, 65129, 65129, 65096, 65096, 65096, 65096, 65096, 65096, 65096, 65096, 65096, 65069, 65069, 65069, 65069, 65069, 65069, 65069, 65069, 65043, 65043, 65043, 65043, 65043, 65043, 65043, 65043, 65043, 65010, 65010, 65010, 65010, 65010, 65010, 65010, 65010, 65010, 64983, 64983, 64983, 64983, 64983, 64983, 64983, 64983, 64950, 64950, 64950, 64950, 64950, 64950, 64950, 64950, 64950, 64924, 64924, 64924, 64924, 64924, 64924, 64924, 64924, 64924, 64891, 64891, 64891, 64891, 64891, 64891, 64891, 64891, 64864, 64864, 64864, 64864, 64864, 64864, 64864, 64864, 64864, 64831, 64831, 64831, 64831, 64831, 64831, 64831, 64831, 64805, 64805, 64805, 64805, 64805, 64805, 64805, 64805, 64805, 64772, 64772, 64772, 64772, 64772, 64772, 64772, 64772, 64746, 64746, 64746, 64746, 64746, 64746, 64746, 64746, 64746, 64713, 64713, 64713, 64713, 64713, 64713, 64713, 64713, 64686, 64686, 64686, 64686, 64686, 64686, 64686, 64686, 64686, 64653, 64653, 64653, 64653, 64653, 64653, 64653, 64653, 64627, 64627, 64627, 64627, 64627, 64627, 64627, 64627, 64627, 64594, 64594, 64594, 64594, 64594, 64594, 64594, 64594, 64568, 64568, 64568, 64568, 64568, 64568, 64568, 64568, 64535, 64535, 64535, 64535, 64535, 64535, 64535, 64535, 64535, 64508, 64508, 64508, 64508, 64508, 64508, 64508, 64508, 64475, 64475, 64475, 64475, 64475, 64475, 64475, 64475, 64449, 64449, 64449, 64449, 64449, 64449, 64449, 64449, 64449, 64416, 64416, 64416, 64416, 64416, 64416, 64416, 64416, 64390, 64390, 64390, 64390, 64390, 64390, 64390, 64390, 64357, 64357, 64357, 64357, 64357, 64357, 64357, 64357, 64357, 64331, 64331, 64331, 64331, 64331, 64331, 64331, 64331, 64298, 64298, 64298, 64298, 64298, 64298, 64298, 64298, 64272, 64272, 64272, 64272, 64272, 64272, 64272, 64272, 64239, 64239, 64239, 64239, 64239, 64239, 64239, 64239, 64239, 64213, 64213, 64213, 64213, 64213, 64213, 64213, 64213, 64180, 64180, 64180, 64180, 64180, 64180, 64180, 64180, 64154, 64154, 64154, 64154, 64154, 64154, 64154, 64154, 64121, 64121, 64121, 64121, 64121, 64121, 64121, 64121, 64095, 64095, 64095, 64095, 64095, 64095, 64095, 64095, 64062, 64062, 64062, 64062, 64062, 64062, 64062, 64062, 64036, 64036, 64036, 64036, 64036, 64036, 64036, 64036, 64036, 64003, 64003, 64003, 64003, 64003, 64003, 64003, 64003, 63977, 63977, 63977, 63977, 63977, 63977, 63977, 63977, 63944, 63944, 63944, 63944, 63944, 63944, 63944, 63944, 63918, 63918, 63918, 63918, 63918, 63918, 63918, 63918, 63886, 63886, 63886, 63886, 63886, 63886, 63886, 63886, 63860, 63860, 63860, 63860, 63860, 63860, 63860, 63860, 63827, 63827, 63827, 63827, 63827, 63827, 63827, 63827, 63801, 63801, 63801, 63801, 63801, 63801, 63801, 63801, 63768, 63768, 63768, 63768, 63768, 63768, 63768, 63768, 63742, 63742, 63742, 63742, 63742, 63742, 63742, 63742, 63716, 63716, 63716, 63716, 63716, 63716, 63716, 63716, 63684, 63684, 63684, 63684, 63684, 63684, 63684, 63684, 63657, 63657, 63657, 63657, 63657, 63657, 63657, 63625, 63625, 63625, 63625, 63625, 63625, 63625, 63625, 63599, 63599, 63599, 63599, 63599, 63599, 63599, 63599, 63566, 63566, 63566, 63566, 63566, 63566, 63566, 63566, 63540, 63540, 63540, 63540, 63540, 63540, 63540, 63540, 63508, 63508, 63508, 63508, 63508, 63508, 63508, 63508, 63482, 63482, 63482, 63482, 63482, 63482, 63482, 63482, 63449, 63449, 63449, 63449, 63449, 63449, 63449, 63423, 63423, 63423, 63423, 63423, 63423, 63423, 63423, 63391, 63391, 63391, 63391, 63391, 63391, 63391, 63391, 63365, 63365, 63365, 63365, 63365, 63365, 63365, 63365, 63332, 63332, 63332, 63332, 63332, 63332, 63332, 63332, 63307, 63307, 63307, 63307, 63307, 63307, 63307, 63274, 63274, 63274, 63274, 63274, 63274, 63274, 63274, 63248, 63248, 63248, 63248, 63248, 63248, 63248, 63248, 63216, 63216, 63216, 63216, 63216, 63216, 63216, 63190, 63190, 63190, 63190, 63190, 63190, 63190, 63190, 63158, 63158, 63158, 63158, 63158, 63158, 63158, 63158, 63132, 63132, 63132, 63132, 63132, 63132, 63132, 63099, 63099, 63099, 63099, 63099, 63099, 63099, 63099, 63073, 63073, 63073, 63073, 63073, 63073, 63073, 63073, 63041, 63041, 63041, 63041, 63041, 63041, 63041, 63015, 63015, 63015, 63015, 63015, 63015, 63015, 63015, 62983, 62983, 62983, 62983, 62983, 62983, 62983, 62983, 62957, 62957, 62957, 62957, 62957, 62957, 62957, 62925, 62925, 62925, 62925, 62925, 62925, 62925, 62925, 62899, 62899, 62899, 62899, 62899, 62899, 62899, 62867, 62867, 62867, 62867, 62867, 62867, 62867, 62867, 62841, 62841, 62841, 62841, 62841, 62841, 62841, 62809, 62809, 62809, 62809, 62809, 62809, 62809, 62809, 62783, 62783, 62783, 62783, 62783, 62783, 62783, 62751, 62751, 62751, 62751, 62751, 62751, 62751, 62751, 62725, 62725, 62725, 62725, 62725, 62725, 62725, 62693, 62693, 62693, 62693, 62693, 62693, 62693, 62693, 62667, 62667, 62667, 62667, 62667, 62667, 62667, 62635, 62635, 62635, 62635, 62635, 62635, 62635, 62635, 62609, 62609, 62609, 62609, 62609, 62609, 62609, 62577, 62577, 62577, 62577, 62577, 62577, 62577, 62577, 62551, 62551, 62551, 62551, 62551, 62551, 62551, 62519, 62519, 62519, 62519, 62519, 62519, 62519, 62519, 62493, 62493, 62493, 62493, 62493, 62493, 62493, 62468, 62468, 62468, 62468, 62468, 62468, 62468, 62436, 62436, 62436, 62436, 62436, 62436, 62436, 62436, 62410, 62410, 62410, 62410, 62410, 62410, 62410, 62378, 62378, 62378, 62378, 62378, 62378, 62378, 62352, 62352, 62352, 62352, 62352, 62352, 62352, 62352, 62320, 62320, 62320, 62320, 62320, 62320, 62320, 62294, 62294, 62294, 62294, 62294, 62294, 62294, 62262, 62262, 62262, 62262, 62262, 62262, 62262, 62262, 62237, 62237, 62237, 62237, 62237, 62237, 62237, 62205, 62205, 62205, 62205, 62205, 62205, 62205, 62179, 62179, 62179, 62179, 62179, 62179, 62179, 62179, 62147, 62147, 62147, 62147, 62147, 62147, 62147, 62122, 62122, 62122, 62122, 62122, 62122, 62122, 62090, 62090, 62090, 62090, 62090, 62090, 62090, 62064, 62064, 62064, 62064, 62064, 62064, 62064, 62064, 62032, 62032, 62032, 62032, 62032, 62032, 62032, 62006, 62006, 62006, 62006, 62006, 62006, 62006, 61975, 61975, 61975, 61975, 61975, 61975, 61975, 61949, 61949, 61949, 61949, 61949, 61949, 61949, 61949, 61917, 61917, 61917, 61917, 61917, 61917, 61917, 61892, 61892, 61892, 61892, 61892, 61892, 61892, 61860, 61860, 61860, 61860, 61860, 61860, 61860, 61834, 61834, 61834, 61834, 61834, 61834, 61834, 61802, 61802, 61802, 61802, 61802, 61802, 61802, 61777, 61777, 61777, 61777, 61777, 61777, 61777, 61745, 61745, 61745, 61745, 61745, 61745, 61745, 61745, 61719, 61719, 61719, 61719, 61719, 61719, 61719, 61688, 61688, 61688, 61688, 61688, 61688, 61688, 61662, 61662, 61662, 61662, 61662, 61662, 61662, 61630, 61630, 61630, 61630, 61630, 61630, 61630, 61605, 61605, 61605, 61605, 61605, 61605, 61605, 61573, 61573, 61573, 61573, 61573, 61573, 61573, 61548, 61548, 61548, 61548, 61548, 61548, 61548, 61516, 61516, 61516, 61516, 61516, 61516, 61516, 61491, 61491, 61491, 61491, 61491, 61491, 61491, 61459, 61459, 61459, 61459, 61459, 61459, 61459, 61433, 61433, 61433, 61433, 61433, 61433, 61433, 61402, 61402, 61402, 61402, 61402, 61402, 61402, 61376, 61376, 61376, 61376, 61376, 61376, 61376, 61345, 61345, 61345, 61345, 61345, 61345, 61345, 61319, 61319, 61319, 61319, 61319, 61319, 61319, 61288, 61288, 61288, 61288, 61288, 61288, 61288, 61262, 61262, 61262, 61262, 61262, 61262, 61262, 61231, 61231, 61231, 61231, 61231, 61231, 61231, 61205, 61205, 61205, 61205, 61205, 61205, 61205, 61180, 61180, 61180, 61180, 61180, 61180, 61180, 61148, 61148, 61148, 61148, 61148, 61148, 61148, 61123, 61123, 61123, 61123, 61123, 61123, 61123, 61091, 61091, 61091, 61091, 61091, 61091, 61091, 61066, 61066, 61066, 61066, 61066, 61066, 61066, 61034, 61034, 61034, 61034, 61034, 61034, 61009, 61009, 61009, 61009, 61009, 61009, 61009, 60978, 60978, 60978, 60978, 60978, 60978, 60978, 60952, 60952, 60952, 60952, 60952, 60952, 60952, 60921, 60921, 60921, 60921, 60921, 60921, 60921, 60896, 60896, 60896, 60896, 60896, 60896, 60896, 60864, 60864, 60864, 60864, 60864, 60864, 60864, 60839, 60839, 60839, 60839, 60839, 60839, 60807, 60807, 60807, 60807, 60807, 60807, 60807, 60782, 60782, 60782, 60782, 60782, 60782, 60782, 60751, 60751, 60751, 60751, 60751, 60751, 60751, 60725, 60725, 60725, 60725, 60725, 60725, 60725, 60694, 60694, 60694, 60694, 60694, 60694, 60669, 60669, 60669, 60669, 60669, 60669, 60669, 60637, 60637, 60637, 60637, 60637, 60637, 60637, 60612, 60612, 60612, 60612, 60612, 60612, 60612, 60581, 60581, 60581, 60581, 60581, 60581, 60556, 60556, 60556, 60556, 60556, 60556, 60556, 60524, 60524, 60524, 60524, 60524, 60524, 60524, 60499, 60499, 60499, 60499, 60499, 60499, 60499, 60468, 60468, 60468, 60468, 60468, 60468, 60442, 60442, 60442, 60442, 60442, 60442, 60442, 60411, 60411, 60411, 60411, 60411, 60411, 60411, 60386, 60386, 60386, 60386, 60386, 60386, 60355, 60355, 60355, 60355, 60355, 60355, 60355, 60330, 60330, 60330, 60330, 60330, 60330, 60330, 60298, 60298, 60298, 60298, 60298, 60298, 60273, 60273, 60273, 60273, 60273, 60273, 60273, 60242, 60242, 60242, 60242, 60242, 60242, 60242, 60217, 60217, 60217, 60217, 60217, 60217, 60185, 60185, 60185, 60185, 60185, 60185, 60185, 60160, 60160, 60160, 60160, 60160, 60160, 60129, 60129, 60129, 60129, 60129, 60129, 60129, 60104, 60104, 60104, 60104, 60104, 60104, 60104, 60073, 60073, 60073, 60073, 60073, 60073, 60048, 60048, 60048, 60048, 60048, 60048, 60048, 60017, 60017, 60017, 60017, 60017, 60017, 59992, 59992, 59992, 59992, 59992, 59992, 59992, 59960, 59960, 59960, 59960, 59960, 59960, 59960, 59935, 59935, 59935, 59935, 59935, 59935, 59910, 59910, 59910, 59910, 59910, 59910, 59910, 59879, 59879, 59879, 59879, 59879, 59879, 59854, 59854, 59854, 59854, 59854, 59854, 59854, 59823, 59823, 59823, 59823, 59823, 59823, 59798, 59798, 59798, 59798, 59798, 59798, 59798, 59767, 59767, 59767, 59767, 59767, 59767, 59742, 59742, 59742, 59742, 59742, 59742, 59742, 59711, 59711, 59711, 59711, 59711, 59711, 59686, 59686, 59686, 59686, 59686, 59686, 59686, 59655, 59655, 59655, 59655, 59655, 59655, 59630, 59630, 59630, 59630, 59630, 59630, 59630, 59599, 59599, 59599, 59599, 59599, 59599, 59574, 59574, 59574, 59574, 59574, 59574, 59574, 59543, 59543, 59543, 59543, 59543, 59543, 59518, 59518, 59518, 59518, 59518, 59518, 59518, 59487, 59487, 59487, 59487, 59487, 59487, 59462, 59462, 59462, 59462, 59462, 59462, 59431, 59431, 59431, 59431, 59431, 59431, 59431, 59406, 59406, 59406, 59406, 59406, 59406, 59375, 59375, 59375, 59375, 59375, 59375, 59375, 59350, 59350, 59350, 59350, 59350, 59350, 59319, 59319, 59319, 59319, 59319, 59319, 59295, 59295, 59295, 59295, 59295, 59295, 59295, 59264, 59264, 59264, 59264, 59264, 59264, 59239, 59239, 59239, 59239, 59239, 59239, 59239, 59208, 59208, 59208, 59208, 59208, 59208, 59183, 59183, 59183, 59183, 59183, 59183, 59152, 59152, 59152, 59152, 59152, 59152, 59152, 59127, 59127, 59127, 59127, 59127, 59127, 59096, 59096, 59096, 59096, 59096, 59096, 59072, 59072, 59072, 59072, 59072, 59072, 59072, 59041, 59041, 59041, 59041, 59041, 59041, 59016, 59016, 59016, 59016, 59016, 59016, 58985, 58985, 58985, 58985, 58985, 58985, 58985, 58960, 58960, 58960, 58960, 58960, 58960, 58929, 58929, 58929, 58929, 58929, 58929, 58905, 58905, 58905, 58905, 58905, 58905, 58905, 58874, 58874, 58874, 58874, 58874, 58874, 58849, 58849, 58849, 58849, 58849, 58849, 58818, 58818, 58818, 58818, 58818, 58818, 58794, 58794, 58794, 58794, 58794, 58794, 58794, 58763, 58763, 58763, 58763, 58763, 58763, 58738, 58738, 58738, 58738, 58738, 58738, 58707, 58707, 58707, 58707, 58707, 58707, 58683, 58683, 58683, 58683, 58683, 58683, 58683, 58658, 58658, 58658, 58658, 58658, 58658, 58627, 58627, 58627, 58627, 58627, 58627, 58603, 58603, 58603, 58603, 58603, 58603, 58572, 58572, 58572, 58572, 58572, 58572, 58547, 58547, 58547, 58547, 58547, 58547, 58547, 58516, 58516, 58516, 58516, 58516, 58516, 58492, 58492, 58492, 58492, 58492, 58492, 58461, 58461, 58461, 58461, 58461, 58461, 58436, 58436, 58436, 58436, 58436, 58436, 58406, 58406, 58406, 58406, 58406, 58406, 58406, 58381, 58381, 58381, 58381, 58381, 58381, 58350, 58350, 58350, 58350, 58350, 58350, 58326, 58326, 58326, 58326, 58326, 58326, 58295, 58295, 58295, 58295, 58295, 58295, 58271, 58271, 58271, 58271, 58271, 58271, 58240, 58240, 58240, 58240, 58240, 58240, 58215, 58215, 58215, 58215, 58215, 58215, 58215, 58185, 58185, 58185, 58185, 58185, 58185, 58160, 58160, 58160, 58160, 58160, 58160, 58130, 58130, 58130, 58130, 58130, 58130, 58105, 58105, 58105, 58105, 58105, 58105, 58075, 58075, 58075, 58075, 58075, 58075, 58050, 58050, 58050, 58050, 58050, 58050, 58019, 58019, 58019, 58019, 58019, 58019, 57995, 57995, 57995, 57995, 57995, 57995, 57964, 57964, 57964, 57964, 57964, 57964, 57940, 57940, 57940, 57940, 57940, 57940, 57940, 57909, 57909, 57909, 57909, 57909, 57909, 57885, 57885, 57885, 57885, 57885, 57885, 57854, 57854, 57854, 57854, 57854, 57854, 57830, 57830, 57830, 57830, 57830, 57830, 57799, 57799, 57799, 57799, 57799, 57799, 57775, 57775, 57775, 57775, 57775, 57775, 57744, 57744, 57744, 57744, 57744, 57744, 57720, 57720, 57720, 57720, 57720, 57720, 57689, 57689, 57689, 57689, 57689, 57689, 57665, 57665, 57665, 57665, 57665, 57665, 57635, 57635, 57635, 57635, 57635, 57635, 57610, 57610, 57610, 57610, 57610, 57610, 57580, 57580, 57580, 57580, 57580, 57580, 57555, 57555, 57555, 57555, 57555, 57555, 57525, 57525, 57525, 57525, 57525, 57525, 57501, 57501, 57501, 57501, 57501, 57501, 57470, 57470, 57470, 57470, 57470, 57470, 57446, 57446, 57446, 57446, 57446, 57446, 57421, 57421, 57421, 57421, 57421, 57421, 57391, 57391, 57391, 57391, 57391, 57391, 57367, 57367, 57367, 57367, 57367, 57367, 57336, 57336, 57336, 57336, 57336, 57312, 57312, 57312, 57312, 57312, 57312, 57282, 57282, 57282, 57282, 57282, 57282, 57257, 57257, 57257, 57257, 57257, 57257, 57227, 57227, 57227, 57227, 57227, 57227, 57203, 57203, 57203, 57203, 57203, 57203, 57172, 57172, 57172, 57172, 57172, 57172, 57148, 57148, 57148, 57148, 57148, 57148, 57118, 57118, 57118, 57118, 57118, 57118, 57093, 57093, 57093, 57093, 57093, 57093, 57063, 57063, 57063, 57063, 57063, 57063, 57039, 57039, 57039, 57039, 57039, 57009, 57009, 57009, 57009, 57009, 57009, 56984, 56984, 56984, 56984, 56984, 56984, 56954, 56954, 56954, 56954, 56954, 56954, 56930, 56930, 56930, 56930, 56930, 56930, 56900, 56900, 56900, 56900, 56900, 56900, 56875, 56875, 56875, 56875, 56875, 56875, 56845, 56845, 56845, 56845, 56845, 56821, 56821, 56821, 56821, 56821, 56821, 56791, 56791, 56791, 56791, 56791, 56791, 56767, 56767, 56767, 56767, 56767, 56767, 56736, 56736, 56736, 56736, 56736, 56736, 56712, 56712, 56712, 56712, 56712, 56712, 56682, 56682, 56682, 56682, 56682, 56658, 56658, 56658, 56658, 56658, 56658, 56628, 56628, 56628, 56628, 56628, 56628, 56603, 56603, 56603, 56603, 56603, 56603, 56573, 56573, 56573, 56573, 56573, 56573, 56549, 56549, 56549, 56549, 56549, 56519, 56519, 56519, 56519, 56519, 56519, 56495, 56495, 56495, 56495, 56495, 56495, 56465, 56465, 56465, 56465, 56465, 56465, 56441, 56441, 56441, 56441, 56441, 56410, 56410, 56410, 56410, 56410, 56410, 56386, 56386, 56386, 56386, 56386, 56386, 56356, 56356, 56356, 56356, 56356, 56356, 56332, 56332, 56332, 56332, 56332, 56302, 56302, 56302, 56302, 56302, 56302, 56278, 56278, 56278, 56278, 56278, 56278, 56254, 56254, 56254, 56254, 56254, 56254, 56224, 56224, 56224, 56224, 56224, 56200, 56200, 56200, 56200, 56200, 56200, 56170, 56170, 56170, 56170, 56170, 56170, 56146, 56146, 56146, 56146, 56146, 56116, 56116, 56116, 56116, 56116, 56116, 56092, 56092, 56092, 56092, 56092, 56092, 56062, 56062, 56062, 56062, 56062, 56062, 56038, 56038, 56038, 56038, 56038, 56008, 56008, 56008, 56008, 56008, 56008, 55984, 55984, 55984, 55984, 55984, 55984, 55954, 55954, 55954, 55954, 55954, 55930, 55930, 55930, 55930, 55930, 55930, 55900, 55900, 55900, 55900, 55900, 55900, 55876, 55876, 55876, 55876, 55876, 55846, 55846, 55846, 55846, 55846, 55846, 55822, 55822, 55822, 55822, 55822, 55822, 55792, 55792, 55792, 55792, 55792, 55768, 55768, 55768, 55768, 55768, 55768, 55738, 55738, 55738, 55738, 55738, 55714, 55714, 55714, 55714, 55714, 55714, 55684, 55684, 55684, 55684, 55684, 55684, 55660, 55660, 55660, 55660, 55660, 55630, 55630, 55630, 55630, 55630, 55630, 55606, 55606, 55606, 55606, 55606, 55606, 55576, 55576, 55576, 55576, 55576, 55552, 55552, 55552, 55552, 55552, 55552, 55523, 55523, 55523, 55523, 55523, 55499, 55499, 55499, 55499, 55499, 55499, 55469, 55469, 55469, 55469, 55469, 55469, 55445, 55445, 55445, 55445, 55445, 55415, 55415, 55415, 55415, 55415, 55415, 55391, 55391, 55391, 55391, 55391, 55361, 55361, 55361, 55361, 55361, 55361, 55338, 55338, 55338, 55338, 55338, 55308, 55308, 55308, 55308, 55308, 55308, 55284, 55284, 55284, 55284, 55284, 55284, 55254, 55254, 55254, 55254, 55254, 55230, 55230, 55230, 55230, 55230, 55230, 55200, 55200, 55200, 55200, 55200, 55177, 55177, 55177, 55177, 55177, 55177, 55147, 55147, 55147, 55147, 55147, 55123, 55123, 55123, 55123, 55123, 55123, 55093, 55093, 55093, 55093, 55093, 55069, 55069, 55069, 55069, 55069, 55069, 55046, 55046, 55046, 55046, 55046, 55016, 55016, 55016, 55016, 55016, 55016, 54992, 54992, 54992, 54992, 54992, 54962, 54962, 54962, 54962, 54962, 54962, 54939, 54939, 54939, 54939, 54939, 54909, 54909, 54909, 54909, 54909, 54909, 54885, 54885, 54885, 54885, 54885, 54855, 54855, 54855, 54855, 54855, 54855, 54832, 54832, 54832, 54832, 54832, 54802, 54802, 54802, 54802, 54802, 54802, 54778, 54778, 54778, 54778, 54778, 54749, 54749, 54749, 54749, 54749, 54749, 54725, 54725, 54725, 54725, 54725, 54695, 54695, 54695, 54695, 54695, 54695, 54671, 54671, 54671, 54671, 54671, 54642, 54642, 54642, 54642, 54642, 54642, 54618, 54618, 54618, 54618, 54618, 54588, 54588, 54588, 54588, 54588, 54565, 54565, 54565, 54565, 54565, 54565, 54535, 54535, 54535, 54535, 54535, 54511, 54511, 54511, 54511, 54511, 54511, 54482, 54482, 54482, 54482, 54482, 54458, 54458, 54458, 54458, 54458, 54458, 54429, 54429, 54429, 54429, 54429, 54405, 54405, 54405, 54405, 54405, 54375, 54375, 54375, 54375, 54375, 54375, 54352, 54352, 54352, 54352, 54352, 54322, 54322, 54322, 54322, 54322, 54322, 54299, 54299, 54299, 54299, 54299, 54269, 54269, 54269, 54269, 54269, 54245, 54245, 54245, 54245, 54245, 54245, 54216, 54216, 54216, 54216, 54216, 54192, 54192, 54192, 54192, 54192, 54192, 54163, 54163, 54163, 54163, 54163, 54139, 54139, 54139, 54139, 54139, 54110, 54110, 54110, 54110, 54110, 54110, 54086, 54086, 54086, 54086, 54086, 54056, 54056, 54056, 54056, 54056, 54033, 54033, 54033, 54033, 54033, 54033, 54003, 54003, 54003, 54003, 54003, 53980, 53980, 53980, 53980, 53980, 53950, 53950, 53950, 53950, 53950, 53950, 53927, 53927, 53927, 53927, 53927, 53897, 53897, 53897, 53897, 53897, 53897, 53874, 53874, 53874, 53874, 53874, 53850, 53850, 53850, 53850, 53850, 53821, 53821, 53821, 53821, 53821, 53821, 53797, 53797, 53797, 53797, 53797, 53768, 53768, 53768, 53768, 53768, 53744, 53744, 53744, 53744, 53744, 53715, 53715, 53715, 53715, 53715, 53715, 53691, 53691, 53691, 53691, 53691, 53662, 53662, 53662, 53662, 53662, 53638, 53638, 53638, 53638, 53638, 53638, 53609, 53609, 53609, 53609, 53609, 53586, 53586, 53586, 53586, 53586, 53556, 53556, 53556, 53556, 53556, 53556, 53533, 53533, 53533, 53533, 53533, 53503, 53503, 53503, 53503, 53503, 53480, 53480, 53480, 53480, 53480, 53451, 53451, 53451, 53451, 53451, 53451, 53427, 53427, 53427, 53427, 53427, 53398, 53398, 53398, 53398, 53398, 53374, 53374, 53374, 53374, 53374, 53345, 53345, 53345, 53345, 53345, 53345, 53322, 53322, 53322, 53322, 53322, 53292, 53292, 53292, 53292, 53292, 53269, 53269, 53269, 53269, 53269, 53240, 53240, 53240, 53240, 53240, 53240, 53216, 53216, 53216, 53216, 53216, 53187, 53187, 53187, 53187, 53187, 53163, 53163, 53163, 53163, 53163, 53134, 53134, 53134, 53134, 53134, 53134, 53111, 53111, 53111, 53111, 53111, 53081, 53081, 53081, 53081, 53081, 53058, 53058, 53058, 53058, 53058, 53029, 53029, 53029, 53029, 53029, 53029, 53005, 53005, 53005, 53005, 53005, 52976, 52976, 52976, 52976, 52976, 52953, 52953, 52953, 52953, 52953, 52924, 52924, 52924, 52924, 52924, 52900, 52900, 52900, 52900, 52900, 52900, 52871, 52871, 52871, 52871, 52871, 52848, 52848, 52848, 52848, 52848, 52819, 52819, 52819, 52819, 52819, 52795, 52795, 52795, 52795, 52795, 52766, 52766, 52766, 52766, 52766, 52743, 52743, 52743, 52743, 52743, 52743, 52713, 52713, 52713, 52713, 52713, 52690, 52690, 52690, 52690, 52690, 52667, 52667, 52667, 52667, 52667, 52638, 52638, 52638, 52638, 52638, 52614, 52614, 52614, 52614, 52614, 52585, 52585, 52585, 52585, 52585, 52585, 52562, 52562, 52562, 52562, 52562, 52533, 52533, 52533, 52533, 52533, 52510, 52510, 52510, 52510, 52510, 52480, 52480, 52480, 52480, 52480, 52457, 52457, 52457, 52457, 52457, 52428, 52428, 52428, 52428, 52428, 52405, 52405, 52405, 52405, 52405, 52405, 52376, 52376, 52376, 52376, 52376, 52352, 52352, 52352, 52352, 52352, 52323, 52323, 52323, 52323, 52323, 52300, 52300, 52300, 52300, 52300, 52271, 52271, 52271, 52271, 52271, 52248, 52248, 52248, 52248, 52248, 52219, 52219, 52219, 52219, 52219, 52195, 52195, 52195, 52195, 52195, 52195, 52166, 52166, 52166, 52166, 52166, 52143, 52143, 52143, 52143, 52143, 52114, 52114, 52114, 52114, 52114, 52091, 52091, 52091, 52091, 52091, 52062, 52062, 52062, 52062, 52062, 52039, 52039, 52039, 52039, 52039, 52010, 52010, 52010, 52010, 52010, 51987, 51987, 51987, 51987, 51987, 51958, 51958, 51958, 51958, 51958, 51934, 51934, 51934, 51934, 51934, 51905, 51905, 51905, 51905, 51905, 51882, 51882, 51882, 51882, 51882, 51853, 51853, 51853, 51853, 51853, 51853, 51830, 51830, 51830, 51830, 51830, 51801, 51801, 51801, 51801, 51801, 51778, 51778, 51778, 51778, 51778, 51749, 51749, 51749, 51749, 51749, 51726, 51726, 51726, 51726, 51726, 51697, 51697, 51697, 51697, 51697, 51674, 51674, 51674, 51674, 51674, 51645, 51645, 51645, 51645, 51645, 51622, 51622, 51622, 51622, 51622, 51593, 51593, 51593, 51593, 51593, 51570, 51570, 51570, 51570, 51570, 51547, 51547, 51547, 51547, 51547, 51518, 51518, 51518, 51518, 51518, 51495, 51495, 51495, 51495, 51495, 51466, 51466, 51466, 51466, 51466, 51443, 51443, 51443, 51443, 51443, 51414, 51414, 51414, 51414, 51414, 51391, 51391, 51391, 51391, 51391, 51362, 51362, 51362, 51362, 51362, 51339, 51339, 51339, 51339, 51339, 51310, 51310, 51310, 51310, 51310, 51287, 51287, 51287, 51287, 51287, 51258, 51258, 51258, 51258, 51258, 51235, 51235, 51235, 51235, 51235, 51206, 51206, 51206, 51206, 51206, 51183, 51183, 51183, 51183, 51183, 51154, 51154, 51154, 51154, 51154, 51131, 51131, 51131, 51131, 51131, 51102, 51102, 51102, 51102, 51102, 51079, 51079, 51079, 51079, 51079, 51050, 51050, 51050, 51050, 51050, 51027, 51027, 51027, 51027, 51027, 50999, 50999, 50999, 50999, 50999, 50976, 50976, 50976, 50976, 50976, 50947, 50947, 50947, 50947, 50947, 50924, 50924, 50924, 50924, 50924, 50895, 50895, 50895, 50895, 50872, 50872, 50872, 50872, 50872, 50843, 50843, 50843, 50843, 50843, 50820, 50820, 50820, 50820, 50820, 50792, 50792, 50792, 50792, 50792, 50769, 50769, 50769, 50769, 50769, 50740, 50740, 50740, 50740, 50740, 50717, 50717, 50717, 50717, 50717, 50688, 50688, 50688, 50688, 50688, 50665, 50665, 50665, 50665, 50665, 50636, 50636, 50636, 50636, 50636, 50613, 50613, 50613, 50613, 50613, 50585, 50585, 50585, 50585, 50585, 50562, 50562, 50562, 50562, 50533, 50533, 50533, 50533, 50533, 50510, 50510, 50510, 50510, 50510, 50482, 50482, 50482, 50482, 50482, 50459, 50459, 50459, 50459, 50459, 50430, 50430, 50430, 50430, 50430, 50407, 50407, 50407, 50407, 50407, 50384, 50384, 50384, 50384, 50384, 50355, 50355, 50355, 50355, 50355, 50332, 50332, 50332, 50332, 50304, 50304, 50304, 50304, 50304, 50281, 50281, 50281, 50281, 50281, 50252, 50252, 50252, 50252, 50252, 50229, 50229, 50229, 50229, 50229, 50201, 50201, 50201, 50201, 50201, 50178, 50178, 50178, 50178, 50178, 50149, 50149, 50149, 50149, 50149, 50126, 50126, 50126, 50126, 50098, 50098, 50098, 50098, 50098, 50075, 50075, 50075, 50075, 50075, 50046, 50046, 50046, 50046, 50046, 50023, 50023, 50023, 50023, 50023, 49995, 49995, 49995, 49995, 49995, 49972, 49972, 49972, 49972, 49943, 49943, 49943, 49943, 49943, 49921, 49921, 49921, 49921, 49921, 49892, 49892, 49892, 49892, 49892, 49869, 49869, 49869, 49869, 49869, 49841, 49841, 49841, 49841, 49841, 49818, 49818, 49818, 49818, 49789, 49789, 49789, 49789, 49789, 49766, 49766, 49766, 49766, 49766, 49738, 49738, 49738, 49738, 49738, 49715, 49715, 49715, 49715, 49715, 49687, 49687, 49687, 49687, 49687, 49664, 49664, 49664, 49664, 49635, 49635, 49635, 49635, 49635, 49612, 49612, 49612, 49612, 49612, 49584, 49584, 49584, 49584, 49584, 49561, 49561, 49561, 49561, 49561, 49533, 49533, 49533, 49533, 49510, 49510, 49510, 49510, 49510, 49481, 49481, 49481, 49481, 49481, 49459, 49459, 49459, 49459, 49459, 49430, 49430, 49430, 49430, 49407, 49407, 49407, 49407, 49407, 49379, 49379, 49379, 49379, 49379, 49356, 49356, 49356, 49356, 49356, 49328, 49328, 49328, 49328, 49328, 49305, 49305, 49305, 49305, 49276, 49276, 49276, 49276, 49276, 49254, 49254, 49254, 49254, 49254, 49231, 49231, 49231, 49231, 49231, 49203, 49203, 49203, 49203, 49180, 49180, 49180, 49180, 49180, 49151, 49151, 49151, 49151, 49151, 49129, 49129, 49129, 49129, 49129, 49100, 49100, 49100, 49100, 49078, 49078, 49078, 49078, 49078, 49049, 49049, 49049, 49049, 49049, 49026, 49026, 49026, 49026, 49026, 48998, 48998, 48998, 48998, 48975, 48975, 48975, 48975, 48975, 48947, 48947, 48947, 48947, 48947, 48924, 48924, 48924, 48924, 48924, 48896, 48896, 48896, 48896, 48873, 48873, 48873, 48873, 48873, 48845, 48845, 48845, 48845, 48845, 48822, 48822, 48822, 48822, 48794, 48794, 48794, 48794, 48794, 48771, 48771, 48771, 48771, 48771, 48743, 48743, 48743, 48743, 48743, 48720, 48720, 48720, 48720, 48692, 48692, 48692, 48692, 48692, 48669, 48669, 48669, 48669, 48669, 48641, 48641, 48641, 48641, 48618, 48618, 48618, 48618, 48618, 48590, 48590, 48590, 48590, 48590, 48567, 48567, 48567, 48567, 48539, 48539, 48539, 48539, 48539, 48516, 48516, 48516, 48516, 48516, 48488, 48488, 48488, 48488, 48488, 48465, 48465, 48465, 48465, 48437, 48437, 48437, 48437, 48437, 48414, 48414, 48414, 48414, 48414, 48386, 48386, 48386, 48386, 48363, 48363, 48363, 48363, 48363, 48335, 48335, 48335, 48335, 48335, 48312, 48312, 48312, 48312, 48284, 48284, 48284, 48284, 48284, 48262, 48262, 48262, 48262, 48262, 48233, 48233, 48233, 48233, 48211, 48211, 48211, 48211, 48211, 48182, 48182, 48182, 48182, 48182, 48160, 48160, 48160, 48160, 48132, 48132, 48132, 48132, 48132, 48109, 48109, 48109, 48109, 48109, 48086, 48086, 48086, 48086, 48058, 48058, 48058, 48058, 48058, 48036, 48036, 48036, 48036, 48007, 48007, 48007, 48007, 48007, 47985, 47985, 47985, 47985, 47985, 47957, 47957, 47957, 47957, 47934, 47934, 47934, 47934, 47934, 47906, 47906, 47906, 47906, 47906, 47883, 47883, 47883, 47883, 47855, 47855, 47855, 47855, 47855, 47833, 47833, 47833, 47833, 47833, 47804, 47804, 47804, 47804, 47782, 47782, 47782, 47782, 47782, 47754, 47754, 47754, 47754, 47731, 47731, 47731, 47731, 47731, 47703, 47703, 47703, 47703, 47703, 47680, 47680, 47680, 47680, 47652, 47652, 47652, 47652, 47652, 47630, 47630, 47630, 47630, 47602, 47602, 47602, 47602, 47602, 47579, 47579, 47579, 47579, 47579, 47551, 47551, 47551, 47551, 47528, 47528, 47528, 47528, 47528, 47500, 47500, 47500, 47500, 47478, 47478, 47478, 47478, 47478, 47450, 47450, 47450, 47450, 47450, 47427, 47427, 47427, 47427, 47399, 47399, 47399, 47399, 47399, 47377, 47377, 47377, 47377, 47348, 47348, 47348, 47348, 47348, 47326, 47326, 47326, 47326, 47298, 47298, 47298, 47298, 47298, 47275, 47275, 47275, 47275, 47275, 47247, 47247, 47247, 47247, 47225, 47225, 47225, 47225, 47225, 47197, 47197, 47197, 47197, 47174, 47174, 47174, 47174, 47174, 47146, 47146, 47146, 47146, 47124, 47124, 47124, 47124, 47124, 47096, 47096, 47096, 47096, 47096, 47073, 47073, 47073, 47073, 47045, 47045, 47045, 47045, 47045, 47023, 47023, 47023, 47023, 46995, 46995, 46995, 46995, 46995, 46972, 46972, 46972, 46972, 46950, 46950, 46950, 46950, 46950, 46922, 46922, 46922, 46922, 46899, 46899, 46899, 46899, 46899, 46871, 46871, 46871, 46871, 46849, 46849, 46849, 46849, 46849, 46821, 46821, 46821, 46821, 46821, 46798, 46798, 46798, 46798, 46770, 46770, 46770, 46770, 46770, 46748, 46748, 46748, 46748, 46720, 46720, 46720, 46720, 46720, 46698, 46698, 46698, 46698, 46670, 46670, 46670, 46670, 46670, 46647, 46647, 46647, 46647, 46619, 46619, 46619, 46619, 46619, 46597, 46597, 46597, 46597, 46569, 46569, 46569, 46569, 46569, 46546, 46546, 46546, 46546, 46518, 46518, 46518, 46518, 46518, 46496, 46496, 46496, 46496, 46468, 46468, 46468, 46468, 46468, 46446, 46446, 46446, 46446, 46418, 46418, 46418, 46418, 46418, 46395, 46395, 46395, 46395, 46367, 46367, 46367, 46367, 46367, 46345, 46345, 46345, 46345, 46317, 46317, 46317, 46317, 46317, 46295, 46295, 46295, 46295, 46267, 46267, 46267, 46267, 46267, 46244, 46244, 46244, 46244, 46216, 46216, 46216, 46216, 46216, 46194, 46194, 46194, 46194, 46166, 46166, 46166, 46166, 46166, 46144, 46144, 46144, 46144, 46116, 46116, 46116, 46116, 46116, 46094, 46094, 46094, 46094, 46066, 46066, 46066, 46066, 46043, 46043, 46043, 46043, 46043, 46015, 46015, 46015, 46015, 45993, 45993, 45993, 45993, 45993, 45965, 45965, 45965, 45965, 45943, 45943, 45943, 45943, 45943, 45915, 45915, 45915, 45915, 45893, 45893, 45893, 45893, 45893, 45870, 45870, 45870, 45870, 45842, 45842, 45842, 45842, 45842, 45820, 45820, 45820, 45820, 45792, 45792, 45792, 45792, 45770, 45770, 45770, 45770, 45770, 45742, 45742, 45742, 45742, 45720, 45720, 45720, 45720, 45720, 45692, 45692, 45692, 45692, 45670, 45670, 45670, 45670, 45670, 45642, 45642, 45642, 45642, 45619, 45619, 45619, 45619, 45592, 45592, 45592, 45592, 45592, 45569, 45569, 45569, 45569, 45541, 45541, 45541, 45541, 45541, 45519, 45519, 45519, 45519, 45491, 45491, 45491, 45491, 45491, 45469, 45469, 45469, 45469, 45441, 45441, 45441, 45441, 45419, 45419, 45419, 45419, 45419, 45391, 45391, 45391, 45391, 45369, 45369, 45369, 45369, 45369, 45341, 45341, 45341, 45341, 45319, 45319, 45319, 45319, 45291, 45291, 45291, 45291, 45291, 45269, 45269, 45269, 45269, 45241, 45241, 45241, 45241, 45241, 45219, 45219, 45219, 45219, 45191, 45191, 45191, 45191, 45169, 45169, 45169, 45169, 45169, 45141, 45141, 45141, 45141, 45119, 45119, 45119, 45119, 45119, 45091, 45091, 45091, 45091, 45069, 45069, 45069, 45069, 45041, 45041, 45041, 45041, 45041, 45019, 45019, 45019, 45019, 44991, 44991, 44991, 44991, 44991, 44969, 44969, 44969, 44969, 44941, 44941, 44941, 44941, 44919, 44919, 44919, 44919, 44919, 44891, 44891, 44891, 44891, 44869, 44869, 44869, 44869, 44841, 44841, 44841, 44841, 44841, 44819, 44819, 44819, 44819, 44791, 44791, 44791, 44791, 44791, 44769, 44769, 44769, 44769, 44747, 44747, 44747, 44747, 44719, 44719, 44719, 44719, 44719, 44697, 44697, 44697, 44697, 44669, 44669, 44669, 44669, 44647, 44647, 44647, 44647, 44647, 44619, 44619, 44619, 44619, 44597, 44597, 44597, 44597, 44569, 44569, 44569, 44569, 44569, 44547, 44547, 44547, 44547, 44519, 44519, 44519, 44519, 44497, 44497, 44497, 44497, 44497, 44469, 44469, 44469, 44469, 44447, 44447, 44447, 44447, 44419, 44419, 44419, 44419, 44419, 44397, 44397, 44397, 44397, 44370, 44370, 44370, 44370, 44347, 44347, 44347, 44347, 44347, 44320, 44320, 44320, 44320, 44298, 44298, 44298, 44298, 44270, 44270, 44270, 44270, 44270, 44248, 44248, 44248, 44248, 44220, 44220, 44220, 44220, 44198, 44198, 44198, 44198, 44198, 44170, 44170, 44170, 44170, 44148, 44148, 44148, 44148, 44120, 44120, 44120, 44120, 44120, 44098, 44098, 44098, 44098, 44071, 44071, 44071, 44071, 44049, 44049, 44049, 44049, 44049, 44021, 44021, 44021, 44021, 43999, 43999, 43999, 43999, 43971, 43971, 43971, 43971, 43971, 43949, 43949, 43949, 43949, 43921, 43921, 43921, 43921, 43899, 43899, 43899, 43899, 43872, 43872, 43872, 43872, 43872, 43849, 43849, 43849, 43849, 43822, 43822, 43822, 43822, 43800, 43800, 43800, 43800, 43800, 43772, 43772, 43772, 43772, 43750, 43750, 43750, 43750, 43722, 43722, 43722, 43722, 43700, 43700, 43700, 43700, 43700, 43673, 43673, 43673, 43673, 43651, 43651, 43651, 43651, 43628, 43628, 43628, 43628, 43628, 43601, 43601, 43601, 43601, 43579, 43579, 43579, 43579, 43551, 43551, 43551, 43551, 43529, 43529, 43529, 43529, 43529, 43501, 43501, 43501, 43501, 43479, 43479, 43479, 43479, 43452, 43452, 43452, 43452, 43430, 43430, 43430, 43430, 43430, 43402, 43402, 43402, 43402, 43380, 43380, 43380, 43380, 43352, 43352, 43352, 43352, 43352, 43330, 43330, 43330, 43330, 43303, 43303, 43303, 43303, 43281, 43281, 43281, 43281, 43253, 43253, 43253, 43253, 43253, 43231, 43231, 43231, 43231, 43204, 43204, 43204, 43204, 43182, 43182, 43182, 43182, 43154, 43154, 43154, 43154, 43154, 43132, 43132, 43132, 43132, 43104, 43104, 43104, 43104, 43082, 43082, 43082, 43082, 43055, 43055, 43055, 43055, 43033, 43033, 43033, 43033, 43033, 43005, 43005, 43005, 43005, 42983, 42983, 42983, 42983, 42956, 42956, 42956, 42956, 42934, 42934, 42934, 42934, 42934, 42906, 42906, 42906, 42906, 42884, 42884, 42884, 42884, 42856, 42856, 42856, 42856, 42834, 42834, 42834, 42834, 42834, 42807, 42807, 42807, 42807, 42785, 42785, 42785, 42785, 42757, 42757, 42757, 42757, 42735, 42735, 42735, 42735, 42708, 42708, 42708, 42708, 42708, 42686, 42686, 42686, 42686, 42658, 42658, 42658, 42658, 42636, 42636, 42636, 42636, 42609, 42609, 42609, 42609, 42587, 42587, 42587, 42587, 42587, 42559, 42559, 42559, 42559, 42537, 42537, 42537, 42537, 42515, 42515, 42515, 42515, 42488, 42488, 42488, 42488, 42466, 42466, 42466, 42466, 42466, 42438, 42438, 42438, 42438, 42416, 42416, 42416, 42416, 42389, 42389, 42389, 42389, 42367, 42367, 42367, 42367, 42339, 42339, 42339, 42339, 42339, 42317, 42317, 42317, 42317, 42290, 42290, 42290, 42290, 42268, 42268, 42268, 42268, 42240, 42240, 42240, 42240, 42218, 42218, 42218, 42218, 42218, 42191, 42191, 42191, 42191, 42169, 42169, 42169, 42169, 42141, 42141, 42141, 42141, 42119, 42119, 42119, 42119, 42092, 42092, 42092, 42092, 42070, 42070, 42070, 42070, 42070, 42042, 42042, 42042, 42042, 42020, 42020, 42020, 42020, 41993, 41993, 41993, 41993, 41971, 41971, 41971, 41971, 41944, 41944, 41944, 41944, 41922, 41922, 41922, 41922, 41922, 41894, 41894, 41894, 41894, 41872, 41872, 41872, 41872, 41845, 41845, 41845, 41845, 41823, 41823, 41823, 41823, 41795, 41795, 41795, 41795, 41773, 41773, 41773, 41773, 41773, 41746, 41746, 41746, 41746, 41724, 41724, 41724, 41724, 41697, 41697, 41697, 41697, 41675, 41675, 41675, 41675, 41647, 41647, 41647, 41647, 41625, 41625, 41625, 41625, 41598, 41598, 41598, 41598, 41598, 41576, 41576, 41576, 41576, 41548, 41548, 41548, 41548, 41527, 41527, 41527, 41527, 41499, 41499, 41499, 41499, 41477, 41477, 41477, 41477, 41455, 41455, 41455, 41455, 41428, 41428, 41428, 41428, 41428, 41406, 41406, 41406, 41406, 41378, 41378, 41378, 41378, 41357, 41357, 41357, 41357, 41329, 41329, 41329, 41329, 41307, 41307, 41307, 41307, 41280, 41280, 41280, 41280, 41258, 41258, 41258, 41258, 41231, 41231, 41231, 41231, 41209, 41209, 41209, 41209, 41209, 41181, 41181, 41181, 41181, 41159, 41159, 41159, 41159, 41132, 41132, 41132, 41132, 41110, 41110, 41110, 41110, 41083, 41083, 41083, 41083, 41061, 41061, 41061, 41061, 41033, 41033, 41033, 41033, 41011, 41011, 41011, 41011, 40984, 40984, 40984, 40984, 40984, 40962, 40962, 40962, 40962, 40935, 40935, 40935, 40935, 40913, 40913, 40913, 40913, 40885, 40885, 40885, 40885, 40864, 40864, 40864, 40864, 40836, 40836, 40836, 40836, 40814, 40814, 40814, 40814, 40787, 40787, 40787, 40787, 40765, 40765, 40765, 40765, 40738, 40738, 40738, 40738, 40738, 40716, 40716, 40716, 40716, 40688, 40688, 40688, 40688, 40667, 40667, 40667, 40667, 40639, 40639, 40639, 40639, 40617, 40617, 40617, 40617, 40590, 40590, 40590, 40590, 40568, 40568, 40568, 40568, 40541, 40541, 40541, 40541, 40519, 40519, 40519, 40519, 40491, 40491, 40491, 40491, 40470, 40470, 40470, 40470, 40442, 40442, 40442, 40442, 40420, 40420, 40420, 40420, 40420, 40393, 40393, 40393, 40393, 40371, 40371, 40371, 40371, 40349, 40349, 40349, 40349, 40322, 40322, 40322, 40322, 40300, 40300, 40300, 40300, 40273, 40273, 40273, 40273, 40251, 40251, 40251, 40251, 40224, 40224, 40224, 40224, 40202, 40202, 40202, 40202, 40174, 40174, 40174, 40174, 40152, 40152, 40152, 40152, 40125, 40125, 40125, 40125, 40103, 40103, 40103, 40103, 40076, 40076, 40076, 40076, 40054, 40054, 40054, 40054, 40027, 40027, 40027, 40027, 40005, 40005, 40005, 40005, 39978, 39978, 39978, 39978, 39956, 39956, 39956, 39956, 39956, 39928, 39928, 39928, 39928, 39907, 39907, 39907, 39907, 39879, 39879, 39879, 39879, 39857, 39857, 39857, 39857, 39830, 39830, 39830, 39830, 39808, 39808, 39808, 39808, 39781, 39781, 39781, 39781, 39759, 39759, 39759, 39759, 39732, 39732, 39732, 39732, 39710, 39710, 39710, 39710, 39683, 39683, 39683, 39683, 39661, 39661, 39661, 39661, 39634, 39634, 39634, 39634, 39612, 39612, 39612, 39612, 39584, 39584, 39584, 39584, 39563, 39563, 39563, 39563, 39535, 39535, 39535, 39535, 39513, 39513, 39513, 39513, 39486, 39486, 39486, 39486, 39464, 39464, 39464, 39464, 39437, 39437, 39437, 39437, 39415, 39415, 39415, 39415, 39388, 39388, 39388, 39388, 39366, 39366, 39366, 39366, 39339, 39339, 39339, 39339, 39317, 39317, 39317, 39317, 39290, 39290, 39290, 39290, 39268, 39268, 39268, 39268, 39246, 39246, 39246, 39246, 39219, 39219, 39219, 39219, 39197, 39197, 39197, 39197, 39170, 39170, 39170, 39170, 39148, 39148, 39148, 39148, 39121, 39121, 39121, 39121, 39099, 39099, 39099, 39099, 39071, 39071, 39071, 39071, 39050, 39050, 39050, 39050, 39022, 39022, 39022, 39022, 39001, 39001, 39001, 39001, 38973, 38973, 38973, 38973, 38951, 38951, 38951, 38951, 38924, 38924, 38924, 38924, 38902, 38902, 38902, 38902, 38875, 38875, 38875, 38875, 38853, 38853, 38853, 38853, 38826, 38826, 38826, 38826, 38804, 38804, 38804, 38804, 38777, 38777, 38777, 38777, 38755, 38755, 38755, 38755, 38728, 38728, 38728, 38728, 38706, 38706, 38706, 38706, 38679, 38679, 38679, 38679, 38657, 38657, 38657, 38657, 38630, 38630, 38630, 38630, 38608, 38608, 38608, 38608, 38581, 38581, 38581, 38581, 38559, 38559, 38559, 38559, 38532, 38532, 38532, 38532, 38510, 38510, 38510, 38483, 38483, 38483, 38483, 38461, 38461, 38461, 38461, 38434, 38434, 38434, 38434, 38412, 38412, 38412, 38412, 38384, 38384, 38384, 38384, 38363, 38363, 38363, 38363, 38335, 38335, 38335, 38335, 38314, 38314, 38314, 38314, 38286, 38286, 38286, 38286, 38265, 38265, 38265, 38265, 38237, 38237, 38237, 38237, 38216, 38216, 38216, 38216, 38188, 38188, 38188, 38188, 38167, 38167, 38167, 38167, 38145, 38145, 38145, 38145, 38118, 38118, 38118, 38118, 38096, 38096, 38096, 38096, 38068, 38068, 38068, 38068, 38047, 38047, 38047, 38019, 38019, 38019, 38019, 37998, 37998, 37998, 37998, 37970, 37970, 37970, 37970, 37949, 37949, 37949, 37949, 37921, 37921, 37921, 37921, 37900, 37900, 37900, 37900, 37872, 37872, 37872, 37872, 37851, 37851, 37851, 37851, 37823, 37823, 37823, 37823, 37802, 37802, 37802, 37802, 37774, 37774, 37774, 37774, 37753, 37753, 37753, 37753, 37725, 37725, 37725, 37725, 37704, 37704, 37704, 37676, 37676, 37676, 37676, 37655, 37655, 37655, 37655, 37627, 37627, 37627, 37627, 37606, 37606, 37606, 37606, 37578, 37578, 37578, 37578, 37557, 37557, 37557, 37557, 37529, 37529, 37529, 37529, 37508, 37508, 37508, 37508, 37480, 37480, 37480, 37480, 37459, 37459, 37459, 37459, 37431, 37431, 37431, 37410, 37410, 37410, 37410, 37382, 37382, 37382, 37382, 37361, 37361, 37361, 37361, 37333, 37333, 37333, 37333, 37312, 37312, 37312, 37312, 37284, 37284, 37284, 37284, 37263, 37263, 37263, 37263, 37235, 37235, 37235, 37235, 37214, 37214, 37214, 37214, 37186, 37186, 37186, 37165, 37165, 37165, 37165, 37137, 37137, 37137, 37137, 37116, 37116, 37116, 37116, 37088, 37088, 37088, 37088, 37067, 37067, 37067, 37067, 37045, 37045, 37045, 37045, 37018, 37018, 37018, 37018, 36996, 36996, 36996, 36969, 36969, 36969, 36969, 36947, 36947, 36947, 36947, 36920, 36920, 36920, 36920, 36898, 36898, 36898, 36898, 36871, 36871, 36871, 36871, 36849, 36849, 36849, 36849, 36822, 36822, 36822, 36822, 36800, 36800, 36800, 36800, 36773, 36773, 36773, 36751, 36751, 36751, 36751, 36724, 36724, 36724, 36724, 36702, 36702, 36702, 36702, 36675, 36675, 36675, 36675, 36653, 36653, 36653, 36653, 36626, 36626, 36626, 36626, 36604, 36604, 36604, 36577, 36577, 36577, 36577, 36555, 36555, 36555, 36555, 36528, 36528, 36528, 36528, 36506, 36506, 36506, 36506, 36479, 36479, 36479, 36479, 36457, 36457, 36457, 36457, 36430, 36430, 36430, 36408, 36408, 36408, 36408, 36381, 36381, 36381, 36381, 36359, 36359, 36359, 36359, 36332, 36332, 36332, 36332, 36310, 36310, 36310, 36310, 36283, 36283, 36283, 36283, 36261, 36261, 36261, 36234, 36234, 36234, 36234, 36212, 36212, 36212, 36212, 36185, 36185, 36185, 36185, 36163, 36163, 36163, 36163, 36136, 36136, 36136, 36136, 36114, 36114, 36114, 36087, 36087, 36087, 36087, 36065, 36065, 36065, 36065, 36038, 36038, 36038, 36038, 36016, 36016, 36016, 36016, 35995, 35995, 35995, 35995, 35967, 35967, 35967, 35946, 35946, 35946, 35946, 35918, 35918, 35918, 35918, 35897, 35897, 35897, 35897, 35869, 35869, 35869, 35869, 35848, 35848, 35848, 35848, 35820, 35820, 35820, 35799, 35799, 35799, 35799, 35771, 35771, 35771, 35771, 35750, 35750, 35750, 35750, 35722, 35722, 35722, 35722, 35701, 35701, 35701, 35701, 35674, 35674, 35674, 35652, 35652, 35652, 35652, 35625, 35625, 35625, 35625, 35603, 35603, 35603, 35603, 35576, 35576, 35576, 35576, 35554, 35554, 35554, 35527, 35527, 35527, 35527, 35505, 35505, 35505, 35505, 35478, 35478, 35478, 35478, 35456, 35456, 35456, 35456, 35429, 35429, 35429, 35407, 35407, 35407, 35407, 35380, 35380, 35380, 35380, 35358, 35358, 35358, 35358, 35331, 35331, 35331, 35331, 35309, 35309, 35309, 35309, 35282, 35282, 35282, 35260, 35260, 35260, 35260, 35233, 35233, 35233, 35233, 35211, 35211, 35211, 35211, 35184, 35184, 35184, 35184, 35162, 35162, 35162, 35135, 35135, 35135, 35135, 35113, 35113, 35113, 35113, 35086, 35086, 35086, 35086, 35064, 35064, 35064, 35037, 35037, 35037, 35037, 35015, 35015, 35015, 35015, 34988, 34988, 34988, 34988, 34966, 34966, 34966, 34966, 34939, 34939, 34939, 34917, 34917, 34917, 34917, 34895, 34895, 34895, 34895, 34868, 34868, 34868, 34868, 34846, 34846, 34846, 34846, 34819, 34819, 34819, 34797, 34797, 34797, 34797, 34770, 34770, 34770, 34770, 34748, 34748, 34748, 34748, 34721, 34721, 34721, 34699, 34699, 34699, 34699, 34672, 34672, 34672, 34672, 34650, 34650, 34650, 34650, 34623, 34623, 34623, 34623, 34601, 34601, 34601, 34574, 34574, 34574, 34574, 34552, 34552, 34552, 34552, 34525, 34525, 34525, 34525, 34503, 34503, 34503, 34476, 34476, 34476, 34476, 34454, 34454, 34454, 34454, 34427, 34427, 34427, 34427, 34405, 34405, 34405, 34378, 34378, 34378, 34378, 34356, 34356, 34356, 34356, 34329, 34329, 34329, 34329, 34307, 34307, 34307, 34280, 34280, 34280, 34280, 34258, 34258, 34258, 34258, 34231, 34231, 34231, 34231, 34209, 34209, 34209, 34182, 34182, 34182, 34182, 34160, 34160, 34160, 34160, 34133, 34133, 34133, 34133, 34111, 34111, 34111, 34084, 34084, 34084, 34084, 34062, 34062, 34062, 34062, 34035, 34035, 34035, 34035, 34013, 34013, 34013, 33986, 33986, 33986, 33986, 33964, 33964, 33964, 33964, 33937, 33937, 33937, 33937, 33915, 33915, 33915, 33888, 33888, 33888, 33888, 33866, 33866, 33866, 33866, 33839, 33839, 33839, 33839, 33817, 33817, 33817, 33795, 33795, 33795, 33795, 33768, 33768, 33768, 33768, 33746, 33746, 33746, 33746, 33719, 33719, 33719, 33697, 33697, 33697, 33697, 33670, 33670, 33670, 33670, 33648, 33648, 33648, 33648, 33621, 33621, 33621, 33599, 33599, 33599, 33599, 33572, 33572, 33572, 33572, 33550, 33550, 33550, 33523, 33523, 33523, 33523, 33501, 33501, 33501, 33501, 33474, 33474, 33474, 33474, 33452, 33452, 33452, 33425, 33425, 33425, 33425, 33403, 33403, 33403, 33403, 33376, 33376, 33376, 33354, 33354, 33354, 33354, 33327, 33327, 33327, 33327, 33305, 33305, 33305, 33305, 33278, 33278, 33278, 33256, 33256, 33256, 33256, 33229, 33229, 33229, 33229, 33207, 33207, 33207, 33179, 33179, 33179, 33179, 33158, 33158, 33158, 33158, 33130, 33130, 33130, 33130, 33109, 33109, 33109, 33081, 33081, 33081, 33081, 33059, 33059, 33059, 33059, 33032, 33032, 33032, 33010, 33010, 33010, 33010, 32983, 32983, 32983, 32983, 32961, 32961, 32961, 32961, 32934, 32934, 32934, 32912, 32912, 32912, 32912, 32885, 32885, 32885, 32885, 32863, 32863, 32863, 32836, 32836, 32836, 32836, 32814, 32814, 32814, 32814, 32787, 32787, 32787, 32765, 32765, 32765, 32765, 32738, 32738, 32738, 32738, 32716, 32716, 32716, 32716, 32694, 32694, 32694, 32667, 32667, 32667, 32667, 32645, 32645, 32645, 32645, 32618, 32618, 32618, 32596, 32596, 32596, 32596, 32568, 32568, 32568, 32568, 32547, 32547, 32547, 32519, 32519, 32519, 32519, 32498, 32498, 32498, 32498, 32470, 32470, 32470, 32448, 32448, 32448, 32448, 32421, 32421, 32421, 32421, 32399, 32399, 32399, 32372, 32372, 32372, 32372, 32350, 32350, 32350, 32350, 32323, 32323, 32323, 32301, 32301, 32301, 32301, 32274, 32274, 32274, 32274, 32252, 32252, 32252, 32225, 32225, 32225, 32225, 32203, 32203, 32203, 32203, 32175, 32175, 32175, 32154, 32154, 32154, 32154, 32126, 32126, 32126, 32126, 32104, 32104, 32104, 32077, 32077, 32077, 32077, 32055, 32055, 32055, 32055, 32028, 32028, 32028, 32006, 32006, 32006, 32006, 31979, 31979, 31979, 31979, 31957, 31957, 31957, 31930, 31930, 31930, 31930, 31908, 31908, 31908, 31908, 31880, 31880, 31880, 31858, 31858, 31858, 31858, 31831, 31831, 31831, 31831, 31809, 31809, 31809, 31782, 31782, 31782, 31782, 31760, 31760, 31760, 31760, 31733, 31733, 31733, 31711, 31711, 31711, 31711, 31684, 31684, 31684, 31684, 31662, 31662, 31662, 31640, 31640, 31640, 31640, 31612, 31612, 31612, 31612, 31591, 31591, 31591, 31563, 31563, 31563, 31563, 31541, 31541, 31541, 31541, 31514, 31514, 31514, 31492, 31492, 31492, 31492, 31465, 31465, 31465, 31465, 31443, 31443, 31443, 31416, 31416, 31416, 31416, 31394, 31394, 31394, 31366, 31366, 31366, 31366, 31344, 31344, 31344, 31344, 31317, 31317, 31317, 31295, 31295, 31295, 31295, 31268, 31268, 31268, 31268, 31246, 31246, 31246, 31219, 31219, 31219, 31219, 31197, 31197, 31197, 31197, 31169, 31169, 31169, 31147, 31147, 31147, 31147, 31120, 31120, 31120, 31098, 31098, 31098, 31098, 31071, 31071, 31071, 31071, 31049, 31049, 31049, 31021, 31021, 31021, 31021, 31000, 31000, 31000, 31000, 30972, 30972, 30972, 30950, 30950, 30950, 30950, 30923, 30923, 30923, 30901, 30901, 30901, 30901, 30874, 30874, 30874, 30874, 30852, 30852, 30852, 30824, 30824, 30824, 30824, 30802, 30802, 30802, 30802, 30775, 30775, 30775, 30753, 30753, 30753, 30753, 30726, 30726, 30726, 30704, 30704, 30704, 30704, 30676, 30676, 30676, 30676, 30654, 30654, 30654, 30627, 30627, 30627, 30627, 30605, 30605, 30605, 30605, 30578, 30578, 30578, 30556, 30556, 30556, 30556, 30534, 30534, 30534, 30506, 30506, 30506, 30506, 30484, 30484, 30484, 30484, 30457, 30457, 30457, 30435, 30435, 30435, 30435, 30408, 30408, 30408, 30386, 30386, 30386, 30386, 30358, 30358, 30358, 30358, 30336, 30336, 30336, 30309, 30309, 30309, 30309, 30287, 30287, 30287, 30260, 30260, 30260, 30260, 30238, 30238, 30238, 30238, 30210, 30210, 30210, 30188, 30188, 30188, 30188, 30161, 30161, 30161, 30139, 30139, 30139, 30139, 30111, 30111, 30111, 30111, 30089, 30089, 30089, 30062, 30062, 30062, 30062, 30040, 30040, 30040, 30012, 30012, 30012, 30012, 29991, 29991, 29991, 29991, 29963, 29963, 29963, 29941, 29941, 29941, 29941, 29914, 29914, 29914, 29892, 29892, 29892, 29892, 29864, 29864, 29864, 29842, 29842, 29842, 29842, 29815, 29815, 29815, 29815, 29793, 29793, 29793, 29765, 29765, 29765, 29765, 29743, 29743, 29743, 29716, 29716, 29716, 29716, 29694, 29694, 29694, 29694, 29666, 29666, 29666, 29644, 29644, 29644, 29644, 29617, 29617, 29617, 29595, 29595, 29595, 29595, 29567, 29567, 29567, 29545, 29545, 29545, 29545, 29518, 29518, 29518, 29518, 29496, 29496, 29496, 29468, 29468, 29468, 29468, 29446, 29446, 29446, 29424, 29424, 29424, 29424, 29397, 29397, 29397, 29375, 29375, 29375, 29375, 29347, 29347, 29347, 29347, 29325, 29325, 29325, 29298, 29298, 29298, 29298, 29276, 29276, 29276, 29248, 29248, 29248, 29248, 29226, 29226, 29226, 29199, 29199, 29199, 29199, 29177, 29177, 29177, 29177, 29149, 29149, 29149, 29127, 29127, 29127, 29127, 29100, 29100, 29100, 29078, 29078, 29078, 29078, 29050, 29050, 29050, 29028, 29028, 29028, 29028, 29000, 29000, 29000, 28978, 28978, 28978, 28978, 28951, 28951, 28951, 28951, 28929, 28929, 28929, 28901, 28901, 28901, 28901, 28879, 28879, 28879, 28852, 28852, 28852, 28852, 28830, 28830, 28830, 28802, 28802, 28802, 28802, 28780, 28780, 28780, 28752, 28752, 28752, 28752, 28730, 28730, 28730, 28730, 28703, 28703, 28703, 28681, 28681, 28681, 28681, 28653, 28653, 28653, 28631, 28631, 28631, 28631, 28603, 28603, 28603, 28581, 28581, 28581, 28581, 28554, 28554, 28554, 28532, 28532, 28532, 28532, 28504, 28504, 28504, 28482, 28482, 28482, 28482, 28454, 28454, 28454, 28454, 28432, 28432, 28432, 28405, 28405, 28405, 28405, 28383, 28383, 28383, 28355, 28355, 28355, 28355, 28333, 28333, 28333, 28311, 28311, 28311, 28311, 28283, 28283, 28283, 28261, 28261, 28261, 28261, 28233, 28233, 28233, 28211, 28211, 28211, 28211, 28184, 28184, 28184, 28162, 28162, 28162, 28162, 28134, 28134, 28134, 28112, 28112, 28112, 28112, 28084, 28084, 28084, 28084, 28062, 28062, 28062, 28034, 28034, 28034, 28034, 28012, 28012, 28012, 27985, 27985, 27985, 27985, 27963, 27963, 27963, 27935, 27935, 27935, 27935, 27913, 27913, 27913, 27885, 27885, 27885, 27885, 27863, 27863, 27863, 27835, 27835, 27835, 27835, 27813, 27813, 27813, 27785, 27785, 27785, 27785, 27763, 27763, 27763, 27736, 27736, 27736, 27736, 27713, 27713, 27713, 27686, 27686, 27686, 27686, 27664, 27664, 27664, 27636, 27636, 27636, 27636, 27614, 27614, 27614, 27586, 27586, 27586, 27586, 27564, 27564, 27564, 27536, 27536, 27536, 27536, 27514, 27514, 27514, 27486, 27486, 27486, 27486, 27464, 27464, 27464, 27436, 27436, 27436, 27436, 27414, 27414, 27414, 27387, 27387, 27387, 27387, 27364, 27364, 27364, 27337, 27337, 27337, 27337, 27314, 27314, 27314, 27287, 27287, 27287, 27287, 27264, 27264, 27264, 27237, 27237, 27237, 27237, 27215, 27215, 27215, 27192, 27192, 27192, 27192, 27165, 27165, 27165, 27142, 27142, 27142, 27142, 27115, 27115, 27115, 27092, 27092, 27092, 27092, 27065, 27065, 27065, 27042, 27042, 27042, 27042, 27015, 27015, 27015, 26992, 26992, 26992, 26992, 26965, 26965, 26965, 26942, 26942, 26942, 26942, 26915, 26915, 26915, 26892, 26892, 26892, 26892, 26865, 26865, 26865, 26842, 26842, 26842, 26842, 26815, 26815, 26815, 26792, 26792, 26792, 26792, 26765, 26765, 26765, 26742, 26742, 26742, 26742, 26715, 26715, 26715, 26692, 26692, 26692, 26692, 26664, 26664, 26664, 26642, 26642, 26642, 26642, 26614, 26614, 26614, 26592, 26592, 26592, 26592, 26564, 26564, 26564, 26542, 26542, 26542, 26542, 26514, 26514, 26514, 26492, 26492, 26492, 26492, 26464, 26464, 26464, 26442, 26442, 26442, 26442, 26414, 26414, 26414, 26392, 26392, 26392, 26392, 26364, 26364, 26364, 26342, 26342, 26342, 26342, 26314, 26314, 26314, 26291, 26291, 26291, 26264, 26264, 26264, 26264, 26241, 26241, 26241, 26213, 26213, 26213, 26213, 26191, 26191, 26191, 26163, 26163, 26163, 26163, 26141, 26141, 26141, 26119, 26119, 26119, 26119, 26091, 26091, 26091, 26068, 26068, 26068, 26068, 26040, 26040, 26040, 26018, 26018, 26018, 26018, 25990, 25990, 25990, 25968, 25968, 25968, 25968, 25940, 25940, 25940, 25918, 25918, 25918, 25890, 25890, 25890, 25890, 25867, 25867, 25867, 25839, 25839, 25839, 25839, 25817, 25817, 25817, 25789, 25789, 25789, 25789, 25767, 25767, 25767, 25739, 25739, 25739, 25739, 25717, 25717, 25717, 25689, 25689, 25689, 25689, 25666, 25666, 25666, 25638, 25638, 25638, 25638, 25616, 25616, 25616, 25588, 25588, 25588, 25566, 25566, 25566, 25566, 25538, 25538, 25538, 25515, 25515, 25515, 25515, 25487, 25487, 25487, 25465, 25465, 25465, 25465, 25437, 25437, 25437, 25414, 25414, 25414, 25414, 25386, 25386, 25386, 25364, 25364, 25364, 25336, 25336, 25336, 25336, 25314, 25314, 25314, 25286, 25286, 25286, 25286, 25263, 25263, 25263, 25235, 25235, 25235, 25235, 25213, 25213, 25213, 25185, 25185, 25185, 25185, 25162, 25162, 25162, 25134, 25134, 25134, 25112, 25112, 25112, 25112, 25084, 25084, 25084, 25061, 25061, 25061, 25061, 25033, 25033, 25033, 25011, 25011, 25011, 25011, 24989, 24989, 24989, 24960, 24960, 24960, 24960, 24938, 24938, 24938, 24910, 24910, 24910, 24887, 24887, 24887, 24887, 24859, 24859, 24859, 24837, 24837, 24837, 24837, 24809, 24809, 24809, 24786, 24786, 24786, 24786, 24758, 24758, 24758, 24736, 24736, 24736, 24708, 24708, 24708, 24708, 24685, 24685, 24685, 24657, 24657, 24657, 24657, 24635, 24635, 24635, 24607, 24607, 24607, 24607, 24584, 24584, 24584, 24556, 24556, 24556, 24533, 24533, 24533, 24533, 24505, 24505, 24505, 24483, 24483, 24483, 24483, 24455, 24455, 24455, 24432, 24432, 24432, 24432, 24404, 24404, 24404, 24381, 24381, 24381, 24353, 24353, 24353, 24353, 24331, 24331, 24331, 24303, 24303, 24303, 24303, 24280, 24280, 24280, 24252, 24252, 24252, 24229, 24229, 24229, 24229, 24201, 24201, 24201, 24179, 24179, 24179, 24179, 24150, 24150, 24150, 24128, 24128, 24128, 24128, 24100, 24100, 24100, 24077, 24077, 24077, 24049, 24049, 24049, 24049, 24026, 24026, 24026, 23998, 23998, 23998, 23998, 23976, 23976, 23976, 23947, 23947, 23947, 23925, 23925, 23925, 23925, 23897, 23897, 23897, 23874, 23874, 23874, 23874, 23851, 23851, 23851, 23823, 23823, 23823, 23801, 23801, 23801, 23801, 23772, 23772, 23772, 23750, 23750, 23750, 23750, 23721, 23721, 23721, 23699, 23699, 23699, 23671, 23671, 23671, 23671, 23648, 23648, 23648, 23620, 23620, 23620, 23620, 23597, 23597, 23597, 23569, 23569, 23569, 23546, 23546, 23546, 23546, 23518, 23518, 23518, 23495, 23495, 23495, 23495, 23467, 23467, 23467, 23444, 23444, 23444, 23416, 23416, 23416, 23416, 23393, 23393, 23393, 23365, 23365, 23365, 23365, 23342, 23342, 23342, 23314, 23314, 23314, 23291, 23291, 23291, 23291, 23263, 23263, 23263, 23240, 23240, 23240, 23240, 23212, 23212, 23212, 23189, 23189, 23189, 23161, 23161, 23161, 23161, 23138, 23138, 23138, 23110, 23110, 23110, 23110, 23087, 23087, 23087, 23059, 23059, 23059, 23036, 23036, 23036, 23036, 23008, 23008, 23008, 22985, 22985, 22985, 22957, 22957, 22957, 22957, 22934, 22934, 22934, 22905, 22905, 22905, 22905, 22883, 22883, 22883, 22854, 22854, 22854, 22832, 22832, 22832, 22832, 22803, 22803, 22803, 22780, 22780, 22780, 22752, 22752, 22752, 22752, 22729, 22729, 22729, 22706, 22706, 22706, 22706, 22678, 22678, 22678, 22655, 22655, 22655, 22627, 22627, 22627, 22627, 22604, 22604, 22604, 22576, 22576, 22576, 22576, 22553, 22553, 22553, 22524, 22524, 22524, 22502, 22502, 22502, 22502, 22473, 22473, 22473, 22450, 22450, 22450, 22422, 22422, 22422, 22422, 22399, 22399, 22399, 22370, 22370, 22370, 22348, 22348, 22348, 22348, 22319, 22319, 22319, 22296, 22296, 22296, 22296, 22268, 22268, 22268, 22245, 22245, 22245, 22216, 22216, 22216, 22216, 22194, 22194, 22194, 22165, 22165, 22165, 22142, 22142, 22142, 22142, 22114, 22114, 22114, 22091, 22091, 22091, 22062, 22062, 22062, 22062, 22039, 22039, 22039, 22011, 22011, 22011, 22011, 21988, 21988, 21988, 21959, 21959, 21959, 21937, 21937, 21937, 21937, 21908, 21908, 21908, 21885, 21885, 21885, 21856, 21856, 21856, 21856, 21834, 21834, 21834, 21805, 21805, 21805, 21782, 21782, 21782, 21782, 21753, 21753, 21753, 21731, 21731, 21731, 21731, 21702, 21702, 21702, 21679, 21679, 21679, 21650, 21650, 21650, 21650, 21627, 21627, 21627, 21604, 21604, 21604, 21576, 21576, 21576, 21576, 21553, 21553, 21553, 21524, 21524, 21524, 21501, 21501, 21501, 21501, 21473, 21473, 21473, 21450, 21450, 21450, 21421, 21421, 21421, 21421, 21398, 21398, 21398, 21369, 21369, 21369, 21346, 21346, 21346, 21346, 21318, 21318, 21318, 21295, 21295, 21295, 21266, 21266, 21266, 21266, 21243, 21243, 21243, 21214, 21214, 21214, 21191, 21191, 21191, 21191, 21162, 21162, 21162, 21139, 21139, 21139, 21111, 21111, 21111, 21111, 21088, 21088, 21088, 21059, 21059, 21059, 21036, 21036, 21036, 21036, 21007, 21007, 21007, 20984, 20984, 20984, 20984, 20955, 20955, 20955, 20932, 20932, 20932, 20904, 20904, 20904, 20904, 20880, 20880, 20880, 20852, 20852, 20852, 20829, 20829, 20829, 20829, 20800, 20800, 20800, 20777, 20777, 20777, 20748, 20748, 20748, 20748, 20725, 20725, 20725, 20696, 20696, 20696, 20673, 20673, 20673, 20644, 20644, 20644, 20644, 20621, 20621, 20621, 20592, 20592, 20592, 20569, 20569, 20569, 20569, 20540, 20540, 20540, 20517, 20517, 20517, 20488, 20488, 20488, 20488, 20465, 20465, 20465, 20442, 20442, 20442, 20413, 20413, 20413, 20413, 20390, 20390, 20390, 20361, 20361, 20361, 20338, 20338, 20338, 20338, 20309, 20309, 20309, 20286, 20286, 20286, 20257, 20257, 20257, 20257, 20234, 20234, 20234, 20205, 20205, 20205, 20182, 20182, 20182, 20182, 20153, 20153, 20153, 20129, 20129, 20129, 20100, 20100, 20100, 20100, 20077, 20077, 20077, 20048, 20048, 20048, 20025, 20025, 20025, 20025, 19996, 19996, 19996, 19973, 19973, 19973, 19944, 19944, 19944, 19921, 19921, 19921, 19921, 19892, 19892, 19892, 19868, 19868, 19868, 19839, 19839, 19839, 19839, 19816, 19816, 19816, 19787, 19787, 19787, 19764, 19764, 19764, 19764, 19735, 19735, 19735, 19712, 19712, 19712, 19682, 19682, 19682, 19682, 19659, 19659, 19659, 19630, 19630, 19630, 19607, 19607, 19607, 19607, 19578, 19578, 19578, 19555, 19555, 19555, 19525, 19525, 19525, 19502, 19502, 19502, 19502, 19473, 19473, 19473, 19450, 19450, 19450, 19421, 19421, 19421, 19421, 19397, 19397, 19397, 19368, 19368, 19368, 19345, 19345, 19345, 19345, 19316, 19316, 19316, 19292, 19292, 19292, 19269, 19269, 19269, 19240, 19240, 19240, 19240, 19217, 19217, 19217, 19187, 19187, 19187, 19164, 19164, 19164, 19164, 19135, 19135, 19135, 19111, 19111, 19111, 19082, 19082, 19082, 19082, 19059, 19059, 19059, 19030, 19030, 19030, 19006, 19006, 19006, 18977, 18977, 18977, 18977, 18954, 18954, 18954, 18924, 18924, 18924, 18901, 18901, 18901, 18901, 18872, 18872, 18872, 18848, 18848, 18848, 18819, 18819, 18819, 18796, 18796, 18796, 18796, 18766, 18766, 18766, 18743, 18743, 18743, 18714, 18714, 18714, 18714, 18690, 18690, 18690, 18661, 18661, 18661, 18637, 18637, 18637, 18608, 18608, 18608, 18608, 18585, 18585, 18585, 18555, 18555, 18555, 18532, 18532, 18532, 18532, 18502, 18502, 18502, 18479, 18479, 18479, 18450, 18450, 18450, 18426, 18426, 18426, 18426, 18397, 18397, 18397, 18373, 18373, 18373, 18344, 18344, 18344, 18344, 18320, 18320, 18320, 18291, 18291, 18291, 18267, 18267, 18267, 18238, 18238, 18238, 18238, 18215, 18215, 18215, 18185, 18185, 18185, 18162, 18162, 18162, 18162, 18132, 18132, 18132, 18109, 18109, 18109, 18085, 18085, 18085, 18056, 18056, 18056, 18056, 18032, 18032, 18032, 18002, 18002, 18002, 17979, 17979, 17979, 17949, 17949, 17949, 17949, 17926, 17926, 17926, 17896, 17896, 17896, 17873, 17873, 17873, 17873, 17843, 17843, 17843, 17820, 17820, 17820, 17790, 17790, 17790, 17766, 17766, 17766, 17766, 17737, 17737, 17737, 17713, 17713, 17713, 17684, 17684, 17684, 17660, 17660, 17660, 17660, 17631, 17631, 17631, 17607, 17607, 17607, 17577, 17577, 17577, 17554, 17554, 17554, 17554, 17524, 17524, 17524, 17500, 17500, 17500, 17471, 17471, 17471, 17471, 17447, 17447, 17447, 17417, 17417, 17417, 17394, 17394, 17394, 17364, 17364, 17364, 17364, 17340, 17340, 17340, 17311, 17311, 17311, 17287, 17287, 17287, 17257, 17257, 17257, 17257, 17234, 17234, 17234, 17204, 17204, 17204, 17180, 17180, 17180, 17151, 17151, 17151, 17151, 17127, 17127, 17127, 17097, 17097, 17097, 17073, 17073, 17073, 17044, 17044, 17044, 17044, 17020, 17020, 17020, 16990, 16990, 16990, 16966, 16966, 16966, 16937, 16937, 16937, 16937, 16913, 16913, 16913, 16889, 16889, 16889, 16859, 16859, 16859, 16835, 16835, 16835, 16835, 16806, 16806, 16806, 16782, 16782, 16782, 16752, 16752, 16752, 16728, 16728, 16728, 16728, 16698, 16698, 16698, 16674, 16674, 16674, 16645, 16645, 16645, 16621, 16621, 16621, 16621, 16591, 16591, 16591, 16567, 16567, 16567, 16537, 16537, 16537, 16513, 16513, 16513, 16513, 16483, 16483, 16483, 16459, 16459, 16459, 16430, 16430, 16430, 16406, 16406, 16406, 16406, 16376, 16376, 16376, 16352, 16352, 16352, 16322, 16322, 16322, 16298, 16298, 16298, 16298, 16268, 16268, 16268, 16244, 16244, 16244, 16214, 16214, 16214, 16190, 16190, 16190, 16190, 16160, 16160, 16160, 16136, 16136, 16136, 16106, 16106, 16106, 16082, 16082, 16082, 16082, 16052, 16052, 16052, 16028, 16028, 16028, 15998, 15998, 15998, 15974, 15974, 15974, 15944, 15944, 15944, 15944, 15920, 15920, 15920, 15890, 15890, 15890, 15866, 15866, 15866, 15836, 15836, 15836, 15836, 15812, 15812, 15812, 15782, 15782, 15782, 15758, 15758, 15758, 15734, 15734, 15734, 15734, 15704, 15704, 15704, 15680, 15680, 15680, 15650, 15650, 15650, 15626, 15626, 15626, 15596, 15596, 15596, 15596, 15571, 15571, 15571, 15541, 15541, 15541, 15517, 15517, 15517, 15487, 15487, 15487, 15487, 15463, 15463, 15463, 15433, 15433, 15433, 15409, 15409, 15409, 15378, 15378, 15378, 15378, 15354, 15354, 15354, 15324, 15324, 15324, 15300, 15300, 15300, 15270, 15270, 15270, 15246, 15246, 15246, 15246, 15215, 15215, 15215, 15191, 15191, 15191, 15161, 15161, 15161, 15137, 15137, 15137, 15137, 15106, 15106, 15106, 15082, 15082, 15082, 15052, 15052, 15052, 15028, 15028, 15028, 14997, 14997, 14997, 14997, 14973, 14973, 14973, 14943, 14943, 14943, 14919, 14919, 14919, 14888, 14888, 14888, 14864, 14864, 14864, 14864, 14834, 14834, 14834, 14809, 14809, 14809, 14779, 14779, 14779, 14755, 14755, 14755, 14755, 14724, 14724, 14724, 14700, 14700, 14700, 14670, 14670, 14670, 14645, 14645, 14645, 14615, 14615, 14615, 14615, 14591, 14591, 14591, 14560, 14560, 14560, 14536, 14536, 14536, 14512, 14512, 14512, 14481, 14481, 14481, 14481, 14457, 14457, 14457, 14426, 14426, 14426, 14402, 14402, 14402, 14371, 14371, 14371, 14371, 14347, 14347, 14347, 14317, 14317, 14317, 14292, 14292, 14292, 14262, 14262, 14262, 14237, 14237, 14237, 14237, 14207, 14207, 14207, 14182, 14182, 14182, 14152, 14152, 14152, 14127, 14127, 14127, 14097, 14097, 14097, 14097, 14072, 14072, 14072, 14042, 14042, 14042, 14017, 14017, 14017, 13987, 13987, 13987, 13962, 13962, 13962, 13962, 13932, 13932, 13932, 13907, 13907, 13907, 13876, 13876, 13876, 13852, 13852, 13852, 13821, 13821, 13821, 13821, 13797, 13797, 13797, 13766, 13766, 13766, 13742, 13742, 13742, 13711, 13711, 13711, 13686, 13686, 13686, 13686, 13656, 13656, 13656, 13631, 13631, 13631, 13600, 13600, 13600, 13576, 13576, 13576, 13545, 13545, 13545, 13545, 13521, 13521, 13521, 13490, 13490, 13490, 13465, 13465, 13465, 13434, 13434, 13434, 13410, 13410, 13410, 13379, 13379, 13379, 13379, 13354, 13354, 13354, 13324, 13324, 13324, 13299, 13299, 13299, 13274, 13274, 13274, 13243, 13243, 13243, 13243, 13219, 13219, 13219, 13188, 13188, 13188, 13163, 13163, 13163, 13132, 13132, 13132, 13108, 13108, 13108, 13108, 13077, 13077, 13077, 13052, 13052, 13052, 13021, 13021, 13021, 12996, 12996, 12996, 12966, 12966, 12966, 12941, 12941, 12941, 12941, 12910, 12910, 12910, 12885, 12885, 12885, 12854, 12854, 12854, 12829, 12829, 12829, 12798, 12798, 12798, 12798, 12774, 12774, 12774, 12743, 12743, 12743, 12718, 12718, 12718, 12687, 12687, 12687, 12662, 12662, 12662, 12631, 12631, 12631, 12631, 12606, 12606, 12606, 12575, 12575, 12575, 12550, 12550, 12550, 12519, 12519, 12519, 12494, 12494, 12494, 12494, 12463, 12463, 12463, 12438, 12438, 12438, 12407, 12407, 12407, 12382, 12382, 12382, 12351, 12351, 12351, 12326, 12326, 12326, 12326, 12295, 12295, 12295, 12270, 12270, 12270, 12239, 12239, 12239, 12214, 12214, 12214, 12183, 12183, 12183, 12158, 12158, 12158, 12158, 12127, 12127, 12127, 12102, 12102, 12102, 12071, 12071, 12071, 12046, 12046, 12046, 12021, 12021, 12021, 12021, 11990, 11990, 11990, 11965, 11965, 11965, 11933, 11933, 11933, 11908, 11908, 11908, 11877, 11877, 11877, 11852, 11852, 11852, 11852, 11821, 11821, 11821, 11796, 11796, 11796, 11764, 11764, 11764, 11739, 11739, 11739, 11708, 11708, 11708, 11683, 11683, 11683, 11683, 11652, 11652, 11652, 11627, 11627, 11627, 11595, 11595, 11595, 11570, 11570, 11570, 11539, 11539, 11539, 11514, 11514, 11514, 11514, 11482, 11482, 11482, 11457, 11457, 11457, 11426, 11426, 11426, 11400, 11400, 11400, 11369, 11369, 11369, 11344, 11344, 11344, 11312, 11312, 11312, 11312, 11287, 11287, 11287, 11256, 11256, 11256, 11231, 11231, 11231, 11199, 11199, 11199, 11174, 11174, 11174, 11142, 11142, 11142, 11142, 11117, 11117, 11117, 11085, 11085, 11085, 11060, 11060, 11060, 11029, 11029, 11029, 11003, 11003, 11003, 10972, 10972, 10972, 10972, 10947, 10947, 10947, 10915, 10915, 10915, 10890, 10890, 10890, 10858, 10858, 10858, 10833, 10833, 10833, 10807, 10807, 10807, 10776, 10776, 10776, 10776, 10750, 10750, 10750, 10719, 10719, 10719, 10693, 10693, 10693, 10662, 10662, 10662, 10636, 10636, 10636, 10605, 10605, 10605, 10579, 10579, 10579, 10579, 10548, 10548, 10548, 10522, 10522, 10522, 10490, 10490, 10490, 10465, 10465, 10465, 10433, 10433, 10433, 10408, 10408, 10408, 10408, 10376, 10376, 10376, 10351, 10351, 10351, 10319, 10319, 10319, 10293, 10293, 10293, 10261, 10261, 10261, 10236, 10236, 10236, 10204, 10204, 10204, 10204, 10179, 10179, 10179, 10147, 10147, 10147, 10121, 10121, 10121, 10089, 10089, 10089, 10064, 10064, 10064, 10032, 10032, 10032, 10006, 10006, 10006, 10006, 9974, 9974, 9974, 9949, 9949, 9949, 9917, 9917, 9917, 9891, 9891, 9891, 9859, 9859, 9859, 9834, 9834, 9834, 9802, 9802, 9802, 9802, 9776, 9776, 9776, 9744, 9744, 9744, 9718, 9718, 9718, 9686, 9686, 9686, 9661, 9661, 9661, 9629, 9629, 9629, 9603, 9603, 9603, 9571, 9571, 9571, 9571, 9545, 9545, 9545, 9520, 9520, 9520, 9487, 9487, 9487, 9462, 9462, 9462, 9430, 9430, 9430, 9404, 9404, 9404, 9372, 9372, 9372, 9372, 9346, 9346, 9346, 9314, 9314, 9314, 9288, 9288, 9288, 9256, 9256, 9256, 9230, 9230, 9230, 9198, 9198, 9198, 9172, 9172, 9172, 9140, 9140, 9140, 9140, 9114, 9114, 9114, 9082, 9082, 9082, 9056, 9056, 9056, 9024, 9024, 9024, 8998, 8998, 8998, 8965, 8965, 8965, 8940, 8940, 8940, 8907, 8907, 8907, 8907, 8881, 8881, 8881, 8849, 8849, 8849, 8823, 8823, 8823, 8791, 8791, 8791, 8765, 8765, 8765, 8732, 8732, 8732, 8706, 8706, 8706, 8674, 8674, 8674, 8674, 8648, 8648, 8648, 8616, 8616, 8616, 8590, 8590, 8590, 8557, 8557, 8557, 8531, 8531, 8531, 8499, 8499, 8499, 8473, 8473, 8473, 8440, 8440, 8440, 8440, 8414, 8414, 8414, 8382, 8382, 8382, 8356, 8356, 8356, 8323, 8323, 8323, 8297, 8297, 8297, 8264, 8264, 8264, 8238, 8238, 8238, 8212, 8212, 8212, 8212, 8180, 8180, 8180, 8153, 8153, 8153, 8121, 8121, 8121, 8095, 8095, 8095, 8062, 8062, 8062, 8036, 8036, 8036, 8003, 8003, 8003, 7977, 7977, 7977, 7944, 7944, 7944, 7944, 7918, 7918, 7918, 7885, 7885, 7885, 7859, 7859, 7859, 7827, 7827, 7827, 7800, 7800, 7800, 7768, 7768, 7768, 7741, 7741, 7741, 7708, 7708, 7708, 7682, 7682, 7682, 7682, 7649, 7649, 7649, 7623, 7623, 7623, 7590, 7590, 7590, 7564, 7564, 7564, 7531, 7531, 7531, 7505, 7505, 7505, 7472, 7472, 7472, 7446, 7446, 7446, 7413, 7413, 7413, 7413, 7386, 7386, 7386, 7353, 7353, 7353, 7327, 7327, 7327, 7294, 7294, 7294, 7268, 7268, 7268, 7235, 7235, 7235, 7208, 7208, 7208, 7175, 7175, 7175, 7149, 7149, 7149, 7149, 7116, 7116, 7116, 7089, 7089, 7089, 7056, 7056, 7056, 7030, 7030, 7030, 6997, 6997, 6997, 6970, 6970, 6970, 6937, 6937, 6937, 6911, 6911, 6911, 6884, 6884, 6884, 6851, 6851, 6851, 6851, 6825, 6825, 6825, 6791, 6791, 6791, 6765, 6765, 6765, 6732, 6732, 6732, 6705, 6705, 6705, 6672, 6672, 6672, 6645, 6645, 6645, 6612, 6612, 6612, 6585, 6585, 6585, 6552, 6552, 6552, 6552, 6525, 6525, 6525, 6492, 6492, 6492, 6466, 6466, 6466, 6432, 6432, 6432, 6406, 6406, 6406, 6372, 6372, 6372, 6346, 6346, 6346, 6312, 6312, 6312, 6285, 6285, 6285, 6252, 6252, 6252, 6252, 6225, 6225, 6225, 6192, 6192, 6192, 6165, 6165, 6165, 6132, 6132, 6132, 6105, 6105, 6105, 6072, 6072, 6072, 6045, 6045, 6045, 6011, 6011, 6011, 5984, 5984, 5984, 5951, 5951, 5951, 5924, 5924, 5924, 5924, 5891, 5891, 5891, 5864, 5864, 5864, 5830, 5830, 5830, 5803, 5803, 5803, 5770, 5770, 5770, 5743, 5743, 5743, 5709, 5709, 5709, 5682, 5682, 5682, 5649, 5649, 5649, 5622, 5622, 5622, 5588, 5588, 5588, 5561, 5561, 5561, 5561, 5534, 5534, 5534, 5500, 5500, 5500, 5473, 5473, 5473, 5440, 5440, 5440, 5413, 5413, 5413, 5379, 5379, 5379, 5352, 5352, 5352, 5318, 5318, 5318, 5291, 5291, 5291, 5257, 5257, 5257, 5230, 5230, 5230, 5196, 5196, 5196, 5196, 5169, 5169, 5169, 5135, 5135, 5135, 5108, 5108, 5108, 5074, 5074, 5074, 5047, 5047, 5047, 5013, 5013, 5013, 4986, 4986, 4986, 4952, 4952, 4952, 4925, 4925, 4925, 4891, 4891, 4891, 4864, 4864, 4864, 4830, 4830, 4830, 4830, 4803, 4803, 4803, 4769, 4769, 4769, 4741, 4741, 4741, 4707, 4707, 4707, 4680, 4680, 4680, 4646, 4646, 4646, 4619, 4619, 4619, 4585, 4585, 4585, 4557, 4557, 4557, 4523, 4523, 4523, 4496, 4496, 4496, 4462, 4462, 4462, 4434, 4434, 4434, 4434, 4400, 4400, 4400, 4373, 4373, 4373, 4339, 4339, 4339, 4311, 4311, 4311, 4277, 4277, 4277, 4250, 4250, 4250, 4222, 4222, 4222, 4188, 4188, 4188, 4161, 4161, 4161, 4126, 4126, 4126, 4099, 4099, 4099, 4064, 4064, 4064, 4037, 4037, 4037, 4003, 4003, 4003, 4003, 3975, 3975, 3975, 3941, 3941, 3941, 3913, 3913, 3913, 3879, 3879, 3879, 3851, 3851, 3851, 3817, 3817, 3817, 3789, 3789, 3789, 3755, 3755, 3755, 3727, 3727, 3727, 3693, 3693, 3693, 3665, 3665, 3665, 3631, 3631, 3631, 3603, 3603, 3603, 3568, 3568, 3568, 3541, 3541, 3541, 3541, 3506, 3506, 3506, 3478, 3478, 3478, 3444, 3444, 3444, 3416, 3416, 3416, 3381, 3381, 3381, 3354, 3354, 3354, 3319, 3319, 3319, 3291, 3291, 3291, 3257, 3257, 3257, 3229, 3229, 3229, 3194, 3194, 3194, 3166, 3166, 3166, 3132, 3132, 3132, 3104, 3104, 3104, 3069, 3069, 3069, 3041, 3041, 3041, 3041, 3006, 3006, 3006, 2978, 2978, 2978, 2944, 2944, 2944, 2916, 2916, 2916, 2881, 2881, 2881, 2853, 2853, 2853, 2825, 2825, 2825, 2790, 2790, 2790, 2762, 2762, 2762, 2727, 2727, 2727, 2699, 2699, 2699, 2664, 2664, 2664, 2636, 2636, 2636, 2601, 2601, 2601, 2573, 2573, 2573, 2538, 2538, 2538, 2510, 2510, 2510, 2475, 2475, 2475, 2475, 2447, 2447, 2447, 2412, 2412, 2412, 2384, 2384, 2384, 2349, 2349, 2349, 2321, 2321, 2321, 2285, 2285, 2285, 2257, 2257, 2257, 2222, 2222, 2222, 2194, 2194, 2194, 2159, 2159, 2159, 2131, 2131, 2131, 2095, 2095, 2095, 2067, 2067, 2067, 2032, 2032, 2032, 2004, 2004, 2004, 1968, 1968, 1968, 1940, 1940, 1940, 1905, 1905, 1905, 1876, 1876, 1876, 1841, 1841, 1841, 1841, 1813, 1813, 1813, 1777, 1777, 1777, 1749, 1749, 1749, 1714, 1714, 1714, 1685, 1685, 1685, 1650, 1650, 1650, 1621, 1621, 1621, 1586, 1586, 1586, 1558, 1558, 1558, 1522, 1522, 1522, 1494, 1494, 1494, 1458, 1458, 1458, 1430, 1430, 1430, 1401, 1401, 1401, 1366, 1366, 1366, 1337, 1337, 1337, 1301, 1301, 1301, 1273, 1273, 1273, 1237, 1237, 1237, 1209, 1209, 1209, 1173, 1173, 1173, 1144, 1144, 1144, 1144, 1109, 1109, 1109, 1080, 1080, 1080, 1044, 1044, 1044, 1016, 1016, 1016, 980, 980, 980, 951, 951, 951, 916, 916, 916, 887, 887, 887, 851, 851, 851, 822, 822, 822, 787, 787, 787, 758, 758, 758, 722, 722, 722, 693, 693, 693, 657, 657, 657, 628, 628, 628, 592, 592, 592, 564, 564, 564, 528, 528, 528, 499, 499, 499, 463, 463, 463, 434, 434, 434, 398, 398, 398, 369, 369, 369, 333, 333, 333, 304, 304, 304, 268, 268, 268, 268, 239, 239, 239, 203, 203, 203, 174, 174, 174, 138, 138, 138, 109, 109, 109, 73, 73, 73, 44, 44, 44, 7, 7, 7, 71978, 71978, 71978, 71949, 71949, 71949, 71913, 71913, 71913, 71884, 71884, 71884, 71848, 71848, 71848, 71819, 71819, 71819, 71783, 71783, 71783, 71754, 71754, 71754, 71718, 71718, 71718, 71689, 71689, 71689, 71653, 71653, 71653, 71624, 71624, 71624, 71588, 71588, 71588, 71559, 71559, 71559, 71523, 71523, 71523, 71494, 71494, 71494, 71458, 71458, 71458, 71429, 71429, 71429, 71393, 71393, 71393, 71364, 71364, 71364, 71328, 71328, 71328, 71300, 71300, 71300, 71264, 71264, 71264, 71235, 71235, 71235, 71199, 71199, 71199, 71170, 71170, 71170, 71135, 71135, 71135, 71106, 71106, 71106, 71106, 71070, 71070, 71070, 71041, 71041, 71041, 71006, 71006, 71006, 70977, 70977, 70977, 70941, 70941, 70941, 70913, 70913, 70913, 70877, 70877, 70877, 70848, 70848, 70848, 70813, 70813, 70813, 70784, 70784, 70784, 70748, 70748, 70748, 70720, 70720, 70720, 70684, 70684, 70684, 70656, 70656, 70656, 70620, 70620, 70620, 70592, 70592, 70592, 70563, 70563, 70563, 70528, 70528, 70528, 70499, 70499, 70499, 70464, 70464, 70464, 70435, 70435, 70435, 70400, 70400, 70400, 70371, 70371, 70371, 70336, 70336, 70336, 70308, 70308, 70308, 70272, 70272, 70272, 70244, 70244, 70244, 70208, 70208, 70208, 70180, 70180, 70180, 70145, 70145, 70145, 70117, 70117, 70117, 70081, 70081, 70081, 70053, 70053, 70053, 70018, 70018, 70018, 69989, 69989, 69989, 69954, 69954, 69954, 69926, 69926, 69926, 69891, 69891, 69891, 69862, 69862, 69862, 69827, 69827, 69827, 69799, 69799, 69799, 69764, 69764, 69764, 69736, 69736, 69736, 69701, 69701, 69701, 69672, 69672, 69672, 69637, 69637, 69637, 69609, 69609, 69609, 69574, 69574, 69574, 69546, 69546, 69546, 69511, 69511, 69511, 69483, 69483, 69483, 69448, 69448, 69448, 69420, 69420, 69420, 69385, 69385, 69385, 69357, 69357, 69357, 69322, 69322, 69322, 69294, 69294, 69294, 69259, 69259, 69259, 69231, 69231, 69231, 69196, 69196, 69196, 69168, 69168, 69168, 69140, 69140, 69140, 69105, 69105, 69105, 69077, 69077, 69077, 69043, 69043, 69043, 69015, 69015, 69015, 68980, 68980, 68980, 68952, 68952, 68952, 68917, 68917, 68917, 68889, 68889, 68889, 68855, 68855, 68855, 68827, 68827, 68827, 68792, 68792, 68792, 68764, 68764, 68764, 68730, 68730, 68730, 68702, 68702, 68702, 68702, 68667, 68667, 68667, 68639, 68639, 68639, 68605, 68605, 68605, 68577, 68577, 68577, 68542, 68542, 68542, 68515, 68515, 68515, 68480, 68480, 68480, 68452, 68452, 68452, 68418, 68418, 68418, 68390, 68390, 68390, 68356, 68356, 68356, 68328, 68328, 68328, 68294, 68294, 68294, 68266, 68266, 68266, 68231, 68231, 68231, 68204, 68204, 68204, 68169, 68169, 68169, 68142, 68142, 68142, 68107, 68107, 68107, 68080, 68080, 68080, 68046, 68046, 68046, 68018, 68018, 68018, 67984, 67984, 67984, 67956, 67956, 67922, 67922, 67922, 67894, 67894, 67894, 67860, 67860, 67860, 67833, 67833, 67833, 67798, 67798, 67798, 67771, 67771, 67771, 67743, 67743, 67743, 67709, 67709, 67709, 67682, 67682, 67682, 67648, 67648, 67648, 67620, 67620, 67620, 67586, 67586, 67586, 67559, 67559, 67559, 67525, 67525, 67525, 67497, 67497, 67497, 67463, 67463, 67463, 67436, 67436, 67436, 67402, 67402, 67402, 67374, 67374, 67374, 67340, 67340, 67340, 67313, 67313, 67313, 67279, 67279, 67279, 67252, 67252, 67252, 67218, 67218, 67218, 67190, 67190, 67190, 67156, 67156, 67156, 67129, 67129, 67129, 67095, 67095, 67095, 67068, 67068, 67068, 67034, 67034, 67034, 67007, 67007, 67007, 66973, 66973, 66973, 66946, 66946, 66946, 66912, 66912, 66912, 66885, 66885, 66885, 66851, 66851, 66851, 66824, 66824, 66824, 66790, 66790, 66790, 66763, 66763, 66763, 66729, 66729, 66729, 66702, 66702, 66702, 66668, 66668, 66668, 66641, 66641, 66641, 66608, 66608, 66608, 66581, 66581, 66581, 66547, 66547, 66547, 66520, 66520, 66520, 66486, 66486, 66486, 66459, 66459, 66459, 66425, 66425, 66425, 66399, 66399, 66399, 66372, 66372, 66372, 66338, 66338, 66338, 66311, 66311, 66311, 66277, 66277, 66277, 66250, 66250, 66250, 66217, 66217, 66217, 66190, 66190, 66190, 66156, 66156, 66156, 66130, 66130, 66130, 66096, 66096, 66096, 66069, 66069, 66069, 66036, 66036, 66036, 66009, 66009, 66009, 65975, 65975, 65975, 65949, 65949, 65949, 65915, 65915, 65915, 65888, 65888, 65888, 65855, 65855, 65855, 65828, 65828, 65828, 65795, 65795, 65795, 65768, 65768, 65768, 65735, 65735, 65735, 65708, 65708, 65708, 65674, 65674, 65674, 65648, 65648, 65648, 65614, 65614, 65614, 65588, 65588, 65588, 65554, 65554, 65554, 65528, 65528, 65494, 65494, 65494, 65468, 65468, 65468, 65435, 65435, 65435, 65408, 65408, 65408, 65375, 65375, 65375, 65348, 65348, 65348, 65315, 65315, 65315, 65288, 65288, 65288, 65255, 65255, 65255, 65229, 65229, 65229, 65195, 65195, 65195, 65169, 65169, 65169, 65136, 65136, 65136, 65109, 65109, 65109, 65076, 65076, 65076, 65050, 65050, 65050, 65023, 65023, 65023, 64990, 64990, 64990, 64964, 64964, 64964, 64930, 64930, 64930, 64904, 64904, 64904, 64871, 64871, 64871, 64845, 64845, 64845, 64812, 64812, 64812, 64785, 64785, 64785, 64752, 64752, 64752, 64726, 64726, 64726, 64693, 64693, 64693, 64666, 64666, 64666, 64633, 64633, 64633, 64607, 64607, 64607, 64574, 64574, 64574, 64548, 64548, 64548, 64515, 64515, 64515, 64489, 64489, 64489, 64456, 64456, 64456, 64429, 64429, 64429, 64397, 64397, 64370, 64370, 64370, 64337, 64337, 64337, 64311, 64311, 64311, 64278, 64278, 64278, 64252, 64252, 64252, 64219, 64219, 64219, 64193, 64193, 64193, 64160, 64160, 64160, 64134, 64134, 64134, 64101, 64101, 64101, 64075, 64075, 64075, 64043, 64043, 64043, 64016, 64016, 64016, 63984, 63984, 63984, 63958, 63958, 63958, 63925, 63925, 63925, 63899, 63899, 63899, 63866, 63866, 63866, 63840, 63840, 63840, 63807, 63807, 63807, 63781, 63781, 63781, 63755, 63755, 63755, 63723, 63723, 63723, 63697, 63697, 63697, 63664, 63664, 63664, 63638, 63638, 63638, 63605, 63605, 63605, 63579, 63579, 63579, 63547, 63547, 63547, 63521, 63521, 63488, 63488, 63488, 63462, 63462, 63462, 63430, 63430, 63430, 63404, 63404, 63404, 63371, 63371, 63371, 63345, 63345, 63345, 63313, 63313, 63313, 63287, 63287, 63287, 63255, 63255, 63255, 63229, 63229, 63229, 63196, 63196, 63196, 63170, 63170, 63170, 63138, 63138, 63138, 63112, 63112, 63112, 63080, 63080, 63080, 63054, 63054, 63054, 63022, 63022, 63022, 62996, 62996, 62996, 62964, 62964, 62964, 62938, 62938, 62938, 62905, 62905, 62905, 62880, 62880, 62880, 62847, 62847, 62847, 62822, 62822, 62822, 62789, 62789, 62764, 62764, 62764, 62731, 62731, 62731, 62706, 62706, 62706, 62673, 62673, 62673, 62648, 62648, 62648, 62615, 62615, 62615, 62590, 62590, 62590, 62558, 62558, 62558, 62532, 62532, 62532, 62500, 62500, 62500, 62474, 62474, 62474, 62448, 62448, 62448, 62416, 62416, 62416, 62391, 62391, 62391, 62359, 62359, 62359, 62333, 62333, 62333, 62301, 62301, 62301, 62275, 62275, 62275, 62243, 62243, 62243, 62218, 62218, 62218, 62186, 62186, 62186, 62160, 62160, 62160, 62128, 62128, 62102, 62102, 62102, 62070, 62070, 62070, 62045, 62045, 62045, 62013, 62013, 62013, 61987, 61987, 61987, 61955, 61955, 61955, 61930, 61930, 61930, 61898, 61898, 61898, 61872, 61872, 61872, 61841, 61841, 61841, 61815, 61815, 61815, 61783, 61783, 61783, 61758, 61758, 61758, 61726, 61726, 61726, 61700, 61700, 61700, 61669, 61669, 61669, 61643, 61643, 61643, 61611, 61611, 61611, 61586, 61586, 61586, 61554, 61554, 61554, 61529, 61529, 61497, 61497, 61497, 61472, 61472, 61472, 61440, 61440, 61440, 61414, 61414, 61414, 61383, 61383, 61383, 61357, 61357, 61357, 61326, 61326, 61326, 61300, 61300, 61300, 61269, 61269, 61269, 61243, 61243, 61243, 61212, 61212, 61212, 61186, 61186, 61186, 61161, 61161, 61161, 61129, 61129, 61129, 61104, 61104, 61104, 61072, 61072, 61072, 61047, 61047, 61047, 61016, 61016, 61016, 60990, 60990, 60959, 60959, 60959, 60933, 60933, 60933, 60902, 60902, 60902, 60877, 60877, 60877, 60845, 60845, 60845, 60820, 60820, 60820, 60788, 60788, 60788, 60763, 60763, 60763, 60732, 60732, 60732, 60707, 60707, 60707, 60675, 60675, 60675, 60650, 60650, 60650, 60618, 60618, 60618, 60593, 60593, 60593, 60562, 60562, 60562, 60537, 60537, 60537, 60505, 60505, 60480, 60480, 60480, 60449, 60449, 60449, 60424, 60424, 60424, 60392, 60392, 60392, 60367, 60367, 60367, 60336, 60336, 60336, 60311, 60311, 60311, 60279, 60279, 60279, 60254, 60254, 60254, 60223, 60223, 60223, 60198, 60198, 60198, 60167, 60167, 60167, 60142, 60142, 60142, 60110, 60110, 60110, 60085, 60085, 60085, 60054, 60054, 60054, 60029, 60029, 59998, 59998, 59998, 59973, 59973, 59973, 59942, 59942, 59942, 59917, 59917, 59917, 59892, 59892, 59892, 59861, 59861, 59861, 59836, 59836, 59836, 59804, 59804, 59804, 59779, 59779, 59779, 59748, 59748, 59748, 59723, 59723, 59723, 59692, 59692, 59692, 59667, 59667, 59667, 59636, 59636, 59636, 59611, 59611, 59611, 59580, 59580, 59555, 59555, 59555, 59524, 59524, 59524, 59499, 59499, 59499, 59468, 59468, 59468, 59443, 59443, 59443, 59412, 59412, 59412, 59388, 59388, 59388, 59357, 59357, 59357, 59332, 59332, 59332, 59301, 59301, 59301, 59276, 59276, 59276, 59245, 59245, 59245, 59220, 59220, 59220, 59189, 59189, 59189, 59164, 59164, 59164, 59133, 59133, 59109, 59109, 59109, 59078, 59078, 59078, 59053, 59053, 59053, 59022, 59022, 59022, 58997, 58997, 58997, 58966, 58966, 58966, 58942, 58942, 58942, 58911, 58911, 58911, 58886, 58886, 58886, 58855, 58855, 58855, 58831, 58831, 58831, 58800, 58800, 58800, 58775, 58775, 58775, 58744, 58744, 58744, 58720, 58720, 58695, 58695, 58695, 58664, 58664, 58664, 58639, 58639, 58639, 58609, 58609, 58609, 58584, 58584, 58584, 58553, 58553, 58553, 58529, 58529, 58529, 58498, 58498, 58498, 58473, 58473, 58473, 58443, 58443, 58443, 58418, 58418, 58418, 58387, 58387, 58387, 58363, 58363, 58363, 58332, 58332, 58307, 58307, 58307, 58277, 58277, 58277, 58252, 58252, 58252, 58222, 58222, 58222, 58197, 58197, 58197, 58166, 58166, 58166, 58142, 58142, 58142, 58111, 58111, 58111, 58087, 58087, 58087, 58056, 58056, 58056, 58032, 58032, 58032, 58001, 58001, 58001, 57977, 57977, 57977, 57946, 57946, 57922, 57922, 57922, 57891, 57891, 57891, 57867, 57867, 57867, 57836, 57836, 57836, 57812, 57812, 57812, 57781, 57781, 57781, 57757, 57757, 57757, 57726, 57726, 57726, 57702, 57702, 57702, 57671, 57671, 57671, 57647, 57647, 57647, 57616, 57616, 57616, 57592, 57592, 57561, 57561, 57561, 57537, 57537, 57537, 57507, 57507, 57507, 57482, 57482, 57482, 57458, 57458, 57458, 57428, 57428, 57428, 57403, 57403, 57403, 57373, 57373, 57373, 57348, 57348, 57348, 57318, 57318, 57318, 57294, 57294, 57294, 57263, 57263, 57263, 57239, 57239, 57209, 57209, 57209, 57184, 57184, 57184, 57154, 57154, 57154, 57130, 57130, 57130, 57100, 57100, 57100, 57075, 57075, 57075, 57045, 57045, 57045, 57021, 57021, 57021, 56990, 56990, 56990, 56966, 56966, 56966, 56936, 56936, 56936, 56912, 56912, 56912, 56881, 56881, 56857, 56857, 56857, 56827, 56827, 56827, 56803, 56803, 56803, 56773, 56773, 56773, 56748, 56748, 56748, 56718, 56718, 56718, 56694, 56694, 56694, 56664, 56664, 56664, 56640, 56640, 56640, 56609, 56609, 56609, 56585, 56585, 56585, 56555, 56555, 56531, 56531, 56531, 56501, 56501, 56501, 56477, 56477, 56477, 56447, 56447, 56447, 56423, 56423, 56423, 56392, 56392, 56392, 56368, 56368, 56368, 56338, 56338, 56338, 56314, 56314, 56314, 56284, 56284, 56284, 56260, 56260, 56260, 56236, 56236, 56206, 56206, 56206, 56182, 56182, 56182, 56152, 56152, 56152, 56128, 56128, 56128, 56098, 56098, 56098, 56074, 56074, 56074, 56044, 56044, 56044, 56020, 56020, 56020, 55990, 55990, 55990, 55966, 55966, 55966, 55936, 55936, 55936, 55912, 55912, 55882, 55882, 55882, 55858, 55858, 55858, 55828, 55828, 55828, 55804, 55804, 55804, 55774, 55774, 55774, 55750, 55750, 55750, 55720, 55720, 55720, 55696, 55696, 55696, 55666, 55666, 55666, 55642, 55642, 55642, 55612, 55612, 55612, 55588, 55588, 55558, 55558, 55558, 55535, 55535, 55535, 55505, 55505, 55505, 55481, 55481, 55481, 55451, 55451, 55451, 55427, 55427, 55427, 55397, 55397, 55397, 55373, 55373, 55373, 55343, 55343, 55343, 55320, 55320, 55320, 55290, 55290, 55266, 55266, 55266, 55236, 55236, 55236, 55212, 55212, 55212, 55183, 55183, 55183, 55159, 55159, 55159, 55129, 55129, 55129, 55105, 55105, 55105, 55075, 55075, 55075, 55052, 55052, 55052, 55028, 55028, 55028, 54998, 54998, 54974, 54974, 54974, 54945, 54945, 54945, 54921, 54921, 54921, 54891, 54891, 54891, 54867, 54867, 54867, 54838, 54838, 54838, 54814, 54814, 54814, 54784, 54784, 54784, 54760, 54760, 54760, 54731, 54731, 54731, 54707, 54707, 54677, 54677, 54677, 54654, 54654, 54654, 54624, 54624, 54624, 54600, 54600, 54600, 54571, 54571, 54571, 54547, 54547, 54547, 54517, 54517, 54517, 54494, 54494, 54494, 54464, 54464, 54464, 54440, 54440, 54440, 54411, 54411, 54387, 54387, 54387, 54358, 54358, 54358, 54334, 54334, 54334, 54304, 54304, 54304, 54281, 54281, 54281, 54251, 54251, 54251, 54228, 54228, 54228, 54198, 54198, 54198, 54174, 54174, 54174, 54145, 54145, 54145, 54121, 54121, 54092, 54092, 54092, 54068, 54068, 54068, 54039, 54039, 54039, 54015, 54015, 54015, 53986, 53986, 53986, 53962, 53962, 53962, 53933, 53933, 53933, 53909, 53909, 53909, 53880, 53880, 53880, 53856, 53856, 53833, 53833, 53833, 53803, 53803, 53803, 53780, 53780, 53780, 53750, 53750, 53750, 53727, 53727, 53727, 53697, 53697, 53697, 53674, 53674, 53674, 53644, 53644, 53644, 53621, 53621, 53621, 53591, 53591, 53568, 53568, 53568, 53539, 53539, 53539, 53515, 53515, 53515, 53486, 53486, 53486, 53462, 53462, 53462, 53433, 53433, 53433, 53410, 53410, 53410, 53380, 53380, 53380, 53357, 53357, 53357, 53327, 53327, 53327, 53304, 53304, 53275, 53275, 53275, 53251, 53251, 53251, 53222, 53222, 53222, 53199, 53199, 53199, 53169, 53169, 53169, 53146, 53146, 53146, 53117, 53117, 53117, 53093, 53093, 53093, 53064, 53064, 53064, 53041, 53041, 53011, 53011, 53011, 52988, 52988, 52988, 52959, 52959, 52959, 52935, 52935, 52935, 52906, 52906, 52906, 52883, 52883, 52883, 52854, 52854, 52854, 52830, 52830, 52830, 52801, 52801, 52801, 52778, 52778, 52748, 52748, 52748, 52725, 52725, 52725, 52702, 52702, 52702, 52673, 52673, 52673, 52649, 52649, 52649, 52620, 52620, 52620, 52597, 52597, 52597, 52568, 52568, 52568, 52544, 52544, 52515, 52515, 52515, 52492, 52492, 52492, 52463, 52463, 52463, 52440, 52440, 52440, 52411, 52411, 52411, 52387, 52387, 52387, 52358, 52358, 52358, 52335, 52335, 52335, 52306, 52306, 52306, 52283, 52283, 52254, 52254, 52254, 52230, 52230, 52230, 52201, 52201, 52201, 52178, 52178, 52178, 52149, 52149, 52149, 52126, 52126, 52126, 52097, 52097, 52097, 52074, 52074, 52074, 52045, 52045, 52045, 52021, 52021, 51992, 51992, 51992, 51969, 51969, 51969, 51940, 51940, 51940, 51917, 51917, 51917, 51888, 51888, 51888, 51865, 51865, 51865, 51836, 51836, 51836, 51813, 51813, 51813, 51784, 51784, 51761, 51761, 51761, 51732, 51732, 51732, 51708, 51708, 51708, 51680, 51680, 51680, 51656, 51656, 51656, 51627, 51627, 51627, 51604, 51604, 51604, 51575, 51575, 51575, 51552, 51552, 51529, 51529, 51529, 51500, 51500, 51500, 51477, 51477, 51477, 51448, 51448, 51448, 51425, 51425, 51425, 51396, 51396, 51396, 51373, 51373, 51373, 51344, 51344, 51344, 51321, 51321, 51321, 51292, 51292, 51269, 51269, 51269, 51241, 51241, 51241, 51218, 51218, 51218, 51189, 51189, 51189, 51166, 51166, 51166, 51137, 51137, 51137, 51114, 51114, 51114, 51085, 51085, 51085, 51062, 51062, 51033, 51033, 51033, 51010, 51010, 51010, 50981, 50981, 50981, 50958, 50958, 50958, 50930, 50930, 50930, 50907, 50907, 50907, 50878, 50878, 50878, 50855, 50855, 50855, 50826, 50826, 50803, 50803, 50803, 50774, 50774, 50774, 50751, 50751, 50751, 50723, 50723, 50723, 50700, 50700, 50700, 50671, 50671, 50671, 50648, 50648, 50648, 50619, 50619, 50619, 50596, 50596, 50568, 50568, 50568, 50545, 50545, 50545, 50516, 50516, 50516, 50493, 50493, 50493, 50464, 50464, 50464, 50441, 50441, 50441, 50413, 50413, 50413, 50390, 50390, 50390, 50367, 50367, 50338, 50338, 50338, 50315, 50315, 50315, 50287, 50287, 50287, 50264, 50264, 50264, 50235, 50235, 50235, 50212, 50212, 50212, 50184, 50184, 50184, 50161, 50161, 50161, 50132, 50132, 50109, 50109, 50109, 50081, 50081, 50081, 50058, 50058, 50058, 50029, 50029, 50029, 50006, 50006, 50006, 49978, 49978, 49978, 49955, 49955, 49955, 49926, 49926, 49926, 49903, 49903, 49875, 49875, 49875, 49852, 49852, 49852, 49824, 49824, 49824, 49801, 49801, 49801, 49772, 49772, 49772, 49749, 49749, 49749, 49721, 49721, 49721, 49698, 49698, 49669, 49669, 49669, 49647, 49647, 49647, 49618, 49618, 49618, 49595, 49595, 49595, 49567, 49567, 49567, 49544, 49544, 49544, 49516, 49516, 49516, 49493, 49493, 49493, 49464, 49464, 49442, 49442, 49442, 49413, 49413, 49413, 49390, 49390, 49390, 49362, 49362, 49362, 49339, 49339, 49339, 49311, 49311, 49311, 49288, 49288, 49288, 49259, 49259, 49259, 49237, 49237, 49214, 49214, 49214, 49185, 49185, 49185, 49163, 49163, 49163, 49134, 49134, 49134, 49112, 49112, 49112, 49083, 49083, 49083, 49060, 49060, 49060, 49032, 49032, 49009, 49009, 49009, 48981, 48981, 48981, 48958, 48958, 48958, 48930, 48930, 48930, 48907, 48907, 48907, 48879, 48879, 48879, 48856, 48856, 48856, 48828, 48828, 48828, 48805, 48805, 48777, 48777, 48777, 48754, 48754, 48754, 48726, 48726, 48726, 48703, 48703, 48703, 48675, 48675, 48675, 48652, 48652, 48652, 48624, 48624, 48624, 48601, 48601, 48573, 48573, 48573, 48550, 48550, 48550, 48522, 48522, 48522, 48499, 48499, 48499, 48471, 48471, 48471, 48448, 48448, 48448, 48420, 48420, 48420, 48397, 48397, 48397, 48369, 48369, 48346, 48346, 48346, 48318, 48318, 48318, 48296, 48296, 48296, 48267, 48267, 48267, 48245, 48245, 48245, 48216, 48216, 48216, 48194, 48194, 48194, 48166, 48166, 48143, 48143, 48143, 48120, 48120, 48120, 48092, 48092, 48092, 48070, 48070, 48070, 48041, 48041, 48041, 48019, 48019, 48019, 47991, 47991, 47991, 47968, 47968, 47940, 47940, 47940, 47917, 47917, 47917, 47889, 47889, 47889, 47866, 47866, 47866, 47838, 47838, 47838, 47816, 47816, 47816, 47788, 47788, 47788, 47765, 47765, 47737, 47737, 47737, 47714, 47714, 47714, 47686, 47686, 47686, 47664, 47664, 47664, 47635, 47635, 47635, 47613, 47613, 47613, 47585, 47585, 47585, 47562, 47562, 47562, 47534, 47534, 47512, 47512, 47512, 47483, 47483, 47483, 47461, 47461, 47461, 47433, 47433, 47433, 47410, 47410, 47410, 47382, 47382, 47382, 47360, 47360, 47360, 47332, 47332, 47309, 47309, 47309, 47281, 47281, 47281, 47259, 47259, 47259, 47230, 47230, 47230, 47208, 47208, 47208, 47180, 47180, 47180, 47157, 47157, 47157, 47129, 47129, 47107, 47107, 47107, 47079, 47079, 47079, 47056, 47056, 47056, 47028, 47028, 47028, 47006, 47006, 47006, 46983, 46983, 46983, 46955, 46955, 46955, 46933, 46933, 46905, 46905, 46905, 46882, 46882, 46882, 46854, 46854, 46854, 46832, 46832, 46832, 46804, 46804, 46804, 46782, 46782, 46782, 46754, 46754, 46754, 46731, 46731, 46703, 46703, 46703, 46681, 46681, 46681, 46653, 46653, 46653, 46630, 46630, 46630, 46602, 46602, 46602, 46580, 46580, 46580, 46552, 46552, 46552, 46530, 46530, 46502, 46502, 46502, 46479, 46479, 46479, 46451, 46451, 46451, 46429, 46429, 46429, 46401, 46401, 46401, 46379, 46379, 46379, 46351, 46351, 46351, 46328, 46328, 46300, 46300, 46300, 46278, 46278, 46278, 46250, 46250, 46250, 46228, 46228, 46228, 46200, 46200, 46200, 46177, 46177, 46177, 46149, 46149, 46149, 46127, 46127, 46099, 46099, 46099, 46077, 46077, 46077, 46049, 46049, 46049, 46027, 46027, 46027, 45999, 45999, 45999, 45976, 45976, 45976, 45948, 45948, 45926, 45926, 45926, 45898, 45898, 45898, 45876, 45876, 45876, 45854, 45854, 45854, 45826, 45826, 45826, 45803, 45803, 45803, 45775, 45775, 45775, 45753, 45753, 45725, 45725, 45725, 45703, 45703, 45703, 45675, 45675, 45675, 45653, 45653, 45653, 45625, 45625, 45625, 45603, 45603, 45603, 45575, 45575, 45575, 45553, 45553, 45525, 45525, 45525, 45502, 45502, 45502, 45475, 45475, 45475, 45452, 45452, 45452, 45425, 45425, 45425, 45402, 45402, 45402, 45374, 45374, 45374, 45352, 45352, 45324, 45324, 45324, 45302, 45302, 45302, 45274, 45274, 45274, 45252, 45252, 45252, 45224, 45224, 45224, 45202, 45202, 45202, 45174, 45174, 45152, 45152, 45152, 45124, 45124, 45124, 45102, 45102, 45102, 45074, 45074, 45074, 45052, 45052, 45052, 45024, 45024, 45024, 45002, 45002, 45002, 44974, 44974, 44952, 44952, 44952, 44924, 44924, 44924, 44902, 44902, 44902, 44874, 44874, 44874, 44852, 44852, 44852, 44824, 44824, 44824, 44802, 44802, 44802, 44774, 44774, 44752, 44752, 44752, 44730, 44730, 44730, 44702, 44702, 44702, 44680, 44680, 44680, 44652, 44652, 44652, 44630, 44630, 44630, 44602, 44602, 44580, 44580, 44580, 44552, 44552, 44552, 44530, 44530, 44530, 44503, 44503, 44503, 44480, 44480, 44480, 44453, 44453, 44453, 44431, 44431, 44431, 44403, 44403, 44381, 44381, 44381, 44353, 44353, 44353, 44331, 44331, 44331, 44303, 44303, 44303, 44281, 44281, 44281, 44253, 44253, 44253, 44231, 44231, 44231, 44204, 44204, 44181, 44181, 44181, 44154, 44154, 44154, 44132, 44132, 44132, 44104, 44104, 44104, 44082, 44082, 44082, 44054, 44054, 44054, 44032, 44032, 44004, 44004, 44004, 43982, 43982, 43982, 43955, 43955, 43955, 43932, 43932, 43932, 43905, 43905, 43905, 43883, 43883, 43883, 43855, 43855, 43855, 43833, 43833, 43805, 43805, 43805, 43783, 43783, 43783, 43756, 43756, 43756, 43733, 43733, 43733, 43706, 43706, 43706, 43684, 43684, 43684, 43656, 43656, 43634, 43634, 43634, 43612, 43612, 43612, 43584, 43584, 43584, 43562, 43562, 43562, 43535, 43535, 43535, 43513, 43513, 43513, 43485, 43485, 43485, 43463, 43463, 43435, 43435, 43435, 43413, 43413, 43413, 43386, 43386, 43386, 43364, 43364, 43364, 43336, 43336, 43336, 43314, 43314, 43314, 43286, 43286, 43264, 43264, 43264, 43237, 43237, 43237, 43215, 43215, 43215, 43187, 43187, 43187, 43165, 43165, 43165, 43137, 43137, 43137, 43115, 43115, 43088, 43088, 43088, 43066, 43066, 43066, 43038, 43038, 43038, 43016, 43016, 43016, 42989, 42989, 42989, 42967, 42967, 42967, 42939, 42939, 42939, 42917, 42917, 42889, 42889, 42889, 42867, 42867, 42867, 42840, 42840, 42840, 42818, 42818, 42818, 42790, 42790, 42790, 42768, 42768, 42768, 42741, 42741, 42719, 42719, 42719, 42691, 42691, 42691, 42669, 42669, 42669, 42642, 42642, 42642, 42620, 42620, 42620, 42592, 42592, 42592, 42570, 42570, 42570, 42548, 42548, 42521, 42521, 42521, 42499, 42499, 42499, 42471, 42471, 42471, 42449, 42449, 42449, 42422, 42422, 42422, 42400, 42400, 42400, 42372, 42372, 42350, 42350, 42350, 42323, 42323, 42323, 42301, 42301, 42301, 42273, 42273, 42273, 42251, 42251, 42251, 42224, 42224, 42224, 42202, 42202, 42174, 42174, 42174, 42152, 42152, 42152, 42125, 42125, 42125, 42103, 42103, 42103, 42075, 42075, 42075, 42053, 42053, 42053, 42026, 42026, 42026, 42004, 42004, 41977, 41977, 41977, 41955, 41955, 41955, 41927, 41927, 41927, 41905, 41905, 41905, 41878, 41878, 41878, 41856, 41856, 41856, 41828, 41828, 41806, 41806, 41806, 41779, 41779, 41779, 41757, 41757, 41757, 41730, 41730, 41730, 41708, 41708, 41708, 41680, 41680, 41680, 41658, 41658, 41631, 41631, 41631, 41609, 41609, 41609, 41581, 41581, 41581, 41559, 41559, 41559, 41532, 41532, 41532, 41510, 41510, 41510, 41483, 41483, 41461, 41461, 41461, 41439, 41439, 41439, 41411, 41411, 41411, 41389, 41389, 41389, 41362, 41362, 41362, 41340, 41340, 41340, 41313, 41313, 41313, 41291, 41291, 41263, 41263, 41263, 41241, 41241, 41241, 41214, 41214, 41214, 41192, 41192, 41192, 41165, 41165, 41165, 41143, 41143, 41143, 41115, 41115, 41094, 41094, 41094, 41066, 41066, 41066, 41044, 41044, 41044, 41017, 41017, 41017, 40995, 40995, 40995, 40968, 40968, 40968, 40946, 40946, 40918, 40918, 40918, 40896, 40896, 40896, 40869, 40869, 40869, 40847, 40847, 40847, 40820, 40820, 40820, 40798, 40798, 40798, 40770, 40770, 40749, 40749, 40749, 40721, 40721, 40721, 40699, 40699, 40699, 40672, 40672, 40672, 40650, 40650, 40650, 40623, 40623, 40623, 40601, 40601, 40574, 40574, 40574, 40552, 40552, 40552, 40524, 40524, 40524, 40502, 40502, 40502, 40475, 40475, 40475, 40453, 40453, 40453, 40426, 40426, 40426, 40404, 40404, 40377, 40377, 40377, 40355, 40355, 40355, 40333, 40333, 40333, 40306, 40306, 40306, 40284, 40284, 40284, 40256, 40256, 40256, 40234, 40234, 40207, 40207, 40207, 40185, 40185, 40185, 40158, 40158, 40158, 40136, 40136, 40136, 40109, 40109, 40109, 40087, 40087, 40087, 40060, 40060, 40038, 40038, 40038, 40010, 40010, 40010, 39989, 39989, 39989, 39961, 39961, 39961, 39939, 39939, 39939, 39912, 39912, 39912, 39890, 39890, 39863, 39863, 39863, 39841, 39841, 39841, 39814, 39814, 39814, 39792, 39792, 39792, 39765, 39765, 39765, 39743, 39743, 39743, 39715, 39715, 39694, 39694, 39694, 39666, 39666, 39666, 39644, 39644, 39644, 39617, 39617, 39617, 39595, 39595, 39595, 39568, 39568, 39568, 39546, 39546, 39519, 39519, 39519, 39497, 39497, 39497, 39470, 39470, 39470, 39448, 39448, 39448, 39421, 39421, 39421, 39399, 39399, 39399, 39372, 39372, 39350, 39350, 39350, 39322, 39322, 39322, 39301, 39301, 39301, 39273, 39273, 39273, 39251, 39251, 39251, 39230, 39230, 39230, 39202, 39202, 39202, 39181, 39181, 39153, 39153, 39153, 39131, 39131, 39131, 39104, 39104, 39104, 39082, 39082, 39082, 39055, 39055, 39055, 39033, 39033, 39033, 39006, 39006, 38984, 38984, 38984, 38957, 38957, 38957, 38935, 38935, 38935, 38908, 38908, 38908, 38886, 38886, 38886, 38859, 38859, 38859, 38837, 38837, 38810, 38810, 38810, 38788, 38788, 38788, 38761, 38761, 38761, 38739, 38739, 38739, 38712, 38712, 38712, 38690, 38690, 38690, 38662, 38662, 38641, 38641, 38641, 38613, 38613, 38613, 38592, 38592, 38592, 38564, 38564, 38564, 38543, 38543, 38543, 38515, 38515, 38515, 38493, 38493, 38466, 38466, 38466, 38444, 38444, 38444, 38417, 38417, 38417, 38395, 38395, 38395, 38368, 38368, 38368, 38346, 38346, 38346, 38319, 38319, 38297, 38297, 38297, 38270, 38270, 38270, 38248, 38248, 38248, 38221, 38221, 38221, 38199, 38199, 38199, 38177, 38177, 38177, 38150, 38150, 38128, 38128, 38128, 38101, 38101, 38101, 38079, 38079, 38079, 38052, 38052, 38052, 38030, 38030, 38030, 38003, 38003, 38003, 37981, 37981, 37954, 37954, 37954, 37932, 37932, 37932, 37905, 37905, 37905, 37883, 37883, 37883, 37856, 37856, 37856, 37834, 37834, 37834, 37807, 37807, 37785, 37785, 37785, 37758, 37758, 37758, 37736, 37736, 37736, 37709, 37709, 37709, 37687, 37687, 37687, 37660, 37660, 37660, 37638, 37638, 37611, 37611, 37611, 37589, 37589, 37589, 37562, 37562, 37562, 37540, 37540, 37540, 37513, 37513, 37513, 37491, 37491, 37491, 37464, 37464, 37442, 37442, 37442, 37415, 37415, 37415, 37393, 37393, 37393, 37366, 37366, 37366, 37344, 37344, 37344, 37317, 37317, 37317, 37295, 37295, 37268, 37268, 37268, 37246, 37246, 37246, 37219, 37219, 37219, 37197, 37197, 37197, 37170, 37170, 37170, 37148, 37148, 37148, 37121, 37121, 37099, 37099, 37099, 37078, 37078, 37078, 37050, 37050, 37050, 37029, 37029, 37029, 37001, 37001, 37001, 36980, 36980, 36980, 36952, 36952, 36931, 36931, 36931, 36903, 36903, 36903, 36882, 36882, 36882, 36854, 36854, 36854, 36833, 36833, 36833, 36805, 36805, 36805, 36784, 36784, 36756, 36756, 36756, 36735, 36735, 36735, 36707, 36707, 36707, 36686, 36686, 36686, 36658, 36658, 36658, 36637, 36637, 36637, 36609, 36609, 36588, 36588, 36588, 36560, 36560, 36560, 36539, 36539, 36539, 36512, 36512, 36512, 36490, 36490, 36490, 36463, 36463, 36463, 36441, 36441, 36414, 36414, 36414, 36392, 36392, 36392, 36365, 36365, 36365, 36343, 36343, 36343, 36316, 36316, 36316, 36294, 36294, 36294, 36267, 36267, 36245, 36245, 36245, 36218, 36218, 36218, 36196, 36196, 36196, 36169, 36169, 36169, 36147, 36147, 36147, 36120, 36120, 36120, 36098, 36098, 36071, 36071, 36071, 36049, 36049, 36049, 36022, 36022, 36022, 36000, 36000, 36000, 35978, 35978, 35978, 35951, 35951, 35951, 35929, 35929, 35929, 35902, 35902, 35880, 35880, 35880, 35853, 35853, 35853, 35831, 35831, 35831, 35804, 35804, 35804, 35782, 35782, 35782, 35755, 35755, 35755, 35733, 35733, 35706, 35706, 35706, 35684, 35684, 35684, 35657, 35657, 35657, 35635, 35635, 35635, 35608, 35608, 35608, 35586, 35586, 35586, 35559, 35559, 35537, 35537, 35537, 35510, 35510, 35510, 35488, 35488, 35488, 35461, 35461, 35461, 35440, 35440, 35440, 35412, 35412, 35412, 35391, 35391, 35363, 35363, 35363, 35342, 35342, 35342, 35314, 35314, 35314, 35293, 35293, 35293, 35265, 35265, 35265, 35244, 35244, 35244, 35216, 35216, 35195, 35195, 35195, 35167, 35167, 35167, 35146, 35146, 35146, 35118, 35118, 35118, 35097, 35097, 35097, 35069, 35069, 35069, 35048, 35048, 35020, 35020, 35020, 34999, 34999, 34999, 34971, 34971, 34971, 34950, 34950, 34950, 34922, 34922, 34922, 34901, 34901, 34901, 34879, 34879, 34852, 34852, 34852, 34830, 34830, 34830, 34803, 34803, 34803, 34781, 34781, 34781, 34754, 34754, 34754, 34732, 34732, 34732, 34705, 34705, 34683, 34683, 34683, 34656, 34656, 34656, 34634, 34634, 34634, 34607, 34607, 34607, 34585, 34585, 34585, 34558, 34558, 34558, 34536, 34536, 34509, 34509, 34509, 34487, 34487, 34487, 34460, 34460, 34460, 34438, 34438, 34438, 34411, 34411, 34411, 34389, 34389, 34389, 34362, 34362, 34340, 34340, 34340, 34313, 34313, 34313, 34291, 34291, 34291, 34264, 34264, 34264, 34242, 34242, 34242, 34215, 34215, 34215, 34193, 34193, 34166, 34166, 34166, 34144, 34144, 34144, 34117, 34117, 34117, 34095, 34095, 34095, 34068, 34068, 34068, 34046, 34046, 34046, 34019, 34019, 33997, 33997, 33997, 33970, 33970, 33970, 33948, 33948, 33948, 33921, 33921, 33921, 33899, 33899, 33899, 33872, 33872, 33872, 33850, 33850, 33823, 33823, 33823, 33801, 33801, 33801, 33779, 33779, 33779, 33752, 33752, 33752, 33730, 33730, 33730, 33703, 33703, 33703, 33681, 33681, 33654, 33654, 33654, 33632, 33632, 33632, 33605, 33605, 33605, 33583, 33583, 33583, 33556, 33556, 33556, 33534, 33534, 33534, 33507, 33507, 33485, 33485, 33485, 33457, 33457, 33457, 33436, 33436, 33436, 33408, 33408, 33408, 33387, 33387, 33387, 33359, 33359, 33359, 33338, 33338, 33310, 33310, 33310, 33288, 33288, 33288, 33261, 33261, 33261, 33239, 33239, 33239, 33212, 33212, 33212, 33190, 33190, 33190, 33163, 33163, 33141, 33141, 33141, 33114, 33114, 33114, 33092, 33092, 33092, 33065, 33065, 33065, 33043, 33043, 33043, 33016, 33016, 33016, 32994, 32994, 32967, 32967, 32967, 32945, 32945, 32945, 32918, 32918, 32918, 32896, 32896, 32896, 32869, 32869, 32869, 32847, 32847, 32847, 32819, 32819, 32798, 32798, 32798, 32770, 32770, 32770, 32749, 32749, 32749, 32727, 32727, 32727, 32699, 32699, 32699, 32678, 32678, 32678, 32650, 32650, 32650, 32628, 32628, 32601, 32601, 32601, 32579, 32579, 32579, 32552, 32552, 32552, 32530, 32530, 32530, 32503, 32503, 32503, 32481, 32481, 32481, 32454, 32454, 32432, 32432, 32432, 32405, 32405, 32405, 32383, 32383, 32383, 32356, 32356, 32356, 32334, 32334, 32334, 32306, 32306, 32306, 32285, 32285, 32257, 32257, 32257, 32235, 32235, 32235, 32208, 32208, 32208, 32186, 32186, 32186, 32159, 32159, 32159, 32137, 32137, 32137, 32110, 32110, 32088, 32088, 32088, 32061, 32061, 32061, 32039, 32039, 32039, 32011, 32011, 32011, 31990, 31990, 31990, 31962, 31962, 31962, 31940, 31940, 31913, 31913, 31913, 31891, 31891, 31891, 31864, 31864, 31864, 31842, 31842, 31842, 31815, 31815, 31815, 31793, 31793, 31793, 31766, 31766, 31744, 31744, 31744, 31716, 31716, 31716, 31694, 31694, 31694, 31667, 31667, 31667, 31645, 31645, 31645, 31623, 31623, 31623, 31596, 31596, 31574, 31574, 31574, 31547, 31547, 31547, 31525, 31525, 31525, 31498, 31498, 31498, 31476, 31476, 31476, 31448, 31448, 31448, 31426, 31426, 31426, 31399, 31399, 31377, 31377, 31377, 31350, 31350, 31350, 31328, 31328, 31328, 31301, 31301, 31301, 31279, 31279, 31279, 31251, 31251, 31251, 31230, 31230, 31202, 31202, 31202, 31180, 31180, 31180, 31153, 31153, 31153, 31131, 31131, 31131, 31104, 31104, 31104, 31082, 31082, 31082, 31054, 31054, 31032, 31032, 31032, 31005, 31005, 31005, 30983, 30983, 30983, 30956, 30956, 30956, 30934, 30934, 30934, 30906, 30906, 30906, 30885, 30885, 30857, 30857, 30857, 30835, 30835, 30835, 30808, 30808, 30808, 30786, 30786, 30786, 30759, 30759, 30759, 30737, 30737, 30737, 30709, 30709, 30687, 30687, 30687, 30660, 30660, 30660, 30638, 30638, 30638, 30611, 30611, 30611, 30589, 30589, 30589, 30561, 30561, 30561, 30539, 30539, 30539, 30517, 30517, 30490, 30490, 30490, 30468, 30468, 30468, 30441, 30441, 30441, 30419, 30419, 30419, 30391, 30391, 30391, 30369, 30369, 30369, 30342, 30342, 30320, 30320, 30320, 30292, 30292, 30292, 30270, 30270, 30270, 30243, 30243, 30243, 30221, 30221, 30221, 30194, 30194, 30194, 30172, 30172, 30144, 30144, 30144, 30122, 30122, 30122, 30095, 30095, 30095, 30073, 30073, 30073, 30045, 30045, 30045, 30023, 30023, 30023, 29996, 29996, 29974, 29974, 29974, 29947, 29947, 29947, 29925, 29925, 29925, 29897, 29897, 29897, 29875, 29875, 29875, 29848, 29848, 29848, 29826, 29826, 29826, 29798, 29798, 29776, 29776, 29776, 29749, 29749, 29749, 29727, 29727, 29727, 29699, 29699, 29699, 29677, 29677, 29677, 29650, 29650, 29650, 29628, 29628, 29600, 29600, 29600, 29578, 29578, 29578, 29551, 29551, 29551, 29529, 29529, 29529, 29501, 29501, 29501, 29479, 29479, 29479, 29452, 29452, 29430, 29430, 29430, 29408, 29408, 29408, 29380, 29380, 29380, 29358, 29358, 29358, 29331, 29331, 29331, 29309, 29309, 29309, 29281, 29281, 29281, 29259, 29259, 29232, 29232, 29232, 29210, 29210, 29210, 29182, 29182, 29182, 29160, 29160, 29160, 29133, 29133, 29133, 29111, 29111, 29111, 29083, 29083, 29061, 29061, 29061, 29033, 29033, 29033, 29011, 29011, 29011, 28984, 28984, 28984, 28962, 28962, 28962, 28934, 28934, 28934, 28912, 28912, 28912, 28885, 28885, 28863, 28863, 28863, 28835, 28835, 28835, 28813, 28813, 28813, 28785, 28785, 28785, 28763, 28763, 28763, 28736, 28736, 28736, 28714, 28714, 28686, 28686, 28686, 28664, 28664, 28664, 28636, 28636, 28636, 28614, 28614, 28614, 28587, 28587, 28587, 28565, 28565, 28565, 28537, 28537, 28515, 28515, 28515, 28487, 28487, 28487, 28465, 28465, 28465, 28438, 28438, 28438, 28416, 28416, 28416, 28388, 28388, 28388, 28366, 28366, 28366, 28344, 28344, 28316, 28316, 28316, 28294, 28294, 28294, 28267, 28267, 28267, 28244, 28244, 28244, 28217, 28217, 28217, 28195, 28195, 28195, 28167, 28167, 28145, 28145, 28145, 28117, 28117, 28117, 28095, 28095, 28095, 28068, 28068, 28068, 28045, 28045, 28045, 28018, 28018, 28018, 27996, 27996, 27996, 27968, 27968, 27946, 27946, 27946, 27918, 27918, 27918, 27896, 27896, 27896, 27868, 27868, 27868, 27846, 27846, 27846, 27819, 27819, 27819, 27796, 27796, 27769, 27769, 27769, 27747, 27747, 27747, 27719, 27719, 27719, 27697, 27697, 27697, 27669, 27669, 27669, 27647, 27647, 27647, 27619, 27619, 27619, 27597, 27597, 27569, 27569, 27569, 27547, 27547, 27547, 27520, 27520, 27520, 27497, 27497, 27497, 27470, 27470, 27470, 27448, 27448, 27448, 27420, 27420, 27420, 27398, 27398, 27370, 27370, 27370, 27348, 27348, 27348, 27320, 27320, 27320, 27298, 27298, 27298, 27270, 27270, 27270, 27248, 27248, 27248, 27226, 27226, 27198, 27198, 27198, 27176, 27176, 27176, 27148, 27148, 27148, 27126, 27126, 27126, 27098, 27098, 27098, 27076, 27076, 27076, 27048, 27048, 27048, 27026, 27026, 26998, 26998, 26998, 26976, 26976, 26976, 26948, 26948, 26948, 26926, 26926, 26926, 26898, 26898, 26898, 26876, 26876, 26876, 26848, 26848, 26848, 26826, 26826, 26798, 26798, 26798, 26776, 26776, 26776, 26748, 26748, 26748, 26726, 26726, 26726, 26698, 26698, 26698, 26676, 26676, 26676, 26648, 26648, 26626, 26626, 26626, 26598, 26598, 26598, 26575, 26575, 26575, 26548, 26548, 26548, 26525, 26525, 26525, 26498, 26498, 26498, 26475, 26475, 26475, 26447, 26447, 26425, 26425, 26425, 26397, 26397, 26397, 26375, 26375, 26375, 26347, 26347, 26347, 26325, 26325, 26325, 26297, 26297, 26297, 26275, 26275, 26275, 26247, 26247, 26225, 26225, 26225, 26197, 26197, 26197, 26174, 26174, 26174, 26146, 26146, 26146, 26124, 26124, 26124, 26102, 26102, 26102, 26074, 26074, 26074, 26052, 26052, 26024, 26024, 26024, 26001, 26001, 26001, 25973, 25973, 25973, 25951, 25951, 25951, 25923, 25923, 25923, 25901, 25901, 25901, 25873, 25873, 25851, 25851, 25851, 25823, 25823, 25823, 25800, 25800, 25800, 25772, 25772, 25772, 25750, 25750, 25750, 25722, 25722, 25722, 25700, 25700, 25700, 25672, 25672, 25649, 25649, 25649, 25621, 25621, 25621, 25599, 25599, 25599, 25571, 25571, 25571, 25549, 25549, 25549, 25521, 25521, 25521, 25498, 25498, 25498, 25470, 25470, 25448, 25448, 25448, 25420, 25420, 25420, 25398, 25398, 25398, 25370, 25370, 25370, 25347, 25347, 25347, 25319, 25319, 25319, 25297, 25297, 25297, 25269, 25269, 25246, 25246, 25246, 25218, 25218, 25218, 25196, 25196, 25196, 25168, 25168, 25168, 25146, 25146, 25146, 25118, 25118, 25118, 25095, 25095, 25095, 25067, 25067, 25045, 25045, 25045, 25017, 25017, 25017, 24994, 24994, 24994, 24972, 24972, 24972, 24944, 24944, 24944, 24921, 24921, 24921, 24893, 24893, 24893, 24871, 24871, 24843, 24843, 24843, 24820, 24820, 24820, 24792, 24792, 24792, 24770, 24770, 24770, 24741, 24741, 24741, 24719, 24719, 24719, 24691, 24691, 24691, 24668, 24668, 24640, 24640, 24640, 24618, 24618, 24618, 24590, 24590, 24590, 24567, 24567, 24567, 24539, 24539, 24539, 24517, 24517, 24517, 24488, 24488, 24488, 24466, 24466, 24438, 24438, 24438, 24415, 24415, 24415, 24387, 24387, 24387, 24365, 24365, 24365, 24336, 24336, 24336, 24314, 24314, 24314, 24286, 24286, 24286, 24263, 24263, 24263, 24235, 24235, 24212, 24212, 24212, 24184, 24184, 24184, 24162, 24162, 24162, 24134, 24134, 24134, 24111, 24111, 24111, 24083, 24083, 24083, 24060, 24060, 24060, 24032, 24032, 24009, 24009, 24009, 23981, 23981, 23981, 23959, 23959, 23959, 23930, 23930, 23930, 23908, 23908, 23908, 23880, 23880, 23880, 23857, 23857, 23857, 23834, 23834, 23806, 23806, 23806, 23784, 23784, 23784, 23755, 23755, 23755, 23733, 23733, 23733, 23704, 23704, 23704, 23682, 23682, 23682, 23654, 23654, 23654, 23631, 23631, 23603, 23603, 23603, 23580, 23580, 23580, 23552, 23552, 23552, 23529, 23529, 23529, 23501, 23501, 23501, 23478, 23478, 23478, 23450, 23450, 23450, 23427, 23427, 23427, 23399, 23399, 23376, 23376, 23376, 23348, 23348, 23348, 23325, 23325, 23325, 23297, 23297, 23297, 23274, 23274, 23274, 23246, 23246, 23246, 23223, 23223, 23223, 23195, 23195, 23172, 23172, 23172, 23144, 23144, 23144, 23121, 23121, 23121, 23093, 23093, 23093, 23070, 23070, 23070, 23042, 23042, 23042, 23019, 23019, 23019, 22991, 22991, 22991, 22968, 22968, 22940, 22940, 22940, 22917, 22917, 22917, 22888, 22888, 22888, 22866, 22866, 22866, 22837, 22837, 22837, 22815, 22815, 22815, 22786, 22786, 22786, 22763, 22763, 22741, 22741, 22741, 22712, 22712, 22712, 22689, 22689, 22689, 22661, 22661, 22661, 22638, 22638, 22638, 22610, 22610, 22610, 22587, 22587, 22587, 22558, 22558, 22558, 22536, 22536, 22507, 22507, 22507, 22484, 22484, 22484, 22456, 22456, 22456, 22433, 22433, 22433, 22405, 22405, 22405, 22382, 22382, 22382, 22353, 22353, 22353, 22331, 22331, 22331, 22302, 22302, 22279, 22279, 22279, 22251, 22251, 22251, 22228, 22228, 22228, 22199, 22199, 22199, 22176, 22176, 22176, 22148, 22148, 22148, 22125, 22125, 22125, 22097, 22097, 22074, 22074, 22074, 22045, 22045, 22045, 22022, 22022, 22022, 21994, 21994, 21994, 21971, 21971, 21971, 21942, 21942, 21942, 21919, 21919, 21919, 21891, 21891, 21891, 21868, 21868, 21839, 21839, 21839, 21816, 21816, 21816, 21788, 21788, 21788, 21765, 21765, 21765, 21736, 21736, 21736, 21713, 21713, 21713, 21685, 21685, 21685, 21662, 21662, 21662, 21633, 21633, 21610, 21610, 21610, 21587, 21587, 21587, 21559, 21559, 21559, 21536, 21536, 21536, 21507, 21507, 21507, 21484, 21484, 21484, 21455, 21455, 21455, 21432, 21432, 21432, 21404, 21404, 21381, 21381, 21381, 21352, 21352, 21352, 21329, 21329, 21329, 21300, 21300, 21300, 21277, 21277, 21277, 21249, 21249, 21249, 21226, 21226, 21226, 21197, 21197, 21197, 21174, 21174, 21145, 21145, 21145, 21122, 21122, 21122, 21093, 21093, 21093, 21070, 21070, 21070, 21042, 21042, 21042, 21019, 21019, 21019, 20990, 20990, 20990, 20967, 20967, 20967, 20938, 20938, 20915, 20915, 20915, 20886, 20886, 20886, 20863, 20863, 20863, 20834, 20834, 20834, 20811, 20811, 20811, 20782, 20782, 20782, 20759, 20759, 20759, 20731, 20731, 20731, 20708, 20708, 20679, 20679, 20679, 20656, 20656, 20656, 20627, 20627, 20627, 20604, 20604, 20604, 20575, 20575, 20575, 20552, 20552, 20552, 20523, 20523, 20523, 20500, 20500, 20500, 20471, 20471, 20471, 20448, 20448, 20425, 20425, 20425, 20396, 20396, 20396, 20373, 20373, 20373, 20344, 20344, 20344, 20320, 20320, 20320, 20292, 20292, 20292, 20268, 20268, 20268, 20239, 20239, 20239, 20216, 20216, 20187, 20187, 20187, 20164, 20164, 20164, 20135, 20135, 20135, 20112, 20112, 20112, 20083, 20083, 20083, 20060, 20060, 20060, 20031, 20031, 20031, 20008, 20008, 20008, 19979, 19979, 19955, 19955, 19955, 19926, 19926, 19926, 19903, 19903, 19903, 19874, 19874, 19874, 19851, 19851, 19851, 19822, 19822, 19822, 19799, 19799, 19799, 19770, 19770, 19770, 19746, 19746, 19746, 19717, 19717, 19694, 19694, 19694, 19665, 19665, 19665, 19642, 19642, 19642, 19613, 19613, 19613, 19589, 19589, 19589, 19560, 19560, 19560, 19537, 19537, 19537, 19508, 19508, 19508, 19485, 19485, 19485, 19456, 19456, 19432, 19432, 19432, 19403, 19403, 19403, 19380, 19380, 19380, 19351, 19351, 19351, 19327, 19327, 19327, 19298, 19298, 19298, 19275, 19275, 19275, 19252, 19252, 19252, 19222, 19222, 19199, 19199, 19199, 19170, 19170, 19170, 19146, 19146, 19146, 19117, 19117, 19117, 19094, 19094, 19094, 19065, 19065, 19065, 19041, 19041, 19041, 19012, 19012, 19012, 18989, 18989, 18989, 18959, 18959, 18936, 18936, 18936, 18907, 18907, 18907, 18883, 18883, 18883, 18854, 18854, 18854, 18831, 18831, 18831, 18801, 18801, 18801, 18778, 18778, 18778, 18749, 18749, 18749, 18725, 18725, 18725, 18696, 18696, 18673, 18673, 18673, 18643, 18643, 18643, 18620, 18620, 18620, 18590, 18590, 18590, 18567, 18567, 18567, 18538, 18538, 18538, 18514, 18514, 18514, 18485, 18485, 18485, 18461, 18461, 18461, 18432, 18432, 18432, 18409, 18409, 18379, 18379, 18379, 18356, 18356, 18356, 18326, 18326, 18326, 18303, 18303, 18303, 18273, 18273, 18273, 18250, 18250, 18250, 18220, 18220, 18220, 18197, 18197, 18197, 18167, 18167, 18167, 18144, 18144, 18120, 18120, 18120, 18091, 18091, 18091, 18067, 18067, 18067, 18038, 18038, 18038, 18014, 18014, 18014, 17985, 17985, 17985, 17961, 17961, 17961, 17932, 17932, 17932, 17908, 17908, 17908, 17879, 17879, 17855, 17855, 17855, 17826, 17826, 17826, 17802, 17802, 17802, 17772, 17772, 17772, 17749, 17749, 17749, 17719, 17719, 17719, 17696, 17696, 17696, 17666, 17666, 17666, 17642, 17642, 17642, 17613, 17613, 17613, 17589, 17589, 17560, 17560, 17560, 17536, 17536, 17536, 17506, 17506, 17506, 17483, 17483, 17483, 17453, 17453, 17453, 17429, 17429, 17429, 17400, 17400, 17400, 17376, 17376, 17376, 17346, 17346, 17346, 17323, 17323, 17323, 17293, 17293, 17269, 17269, 17269, 17240, 17240, 17240, 17216, 17216, 17216, 17186, 17186, 17186, 17162, 17162, 17162, 17133, 17133, 17133, 17109, 17109, 17109, 17079, 17079, 17079, 17055, 17055, 17055, 17026, 17026, 17026, 17002, 17002, 16972, 16972, 16972, 16948, 16948, 16948, 16925, 16925, 16925, 16895, 16895, 16895, 16871, 16871, 16871, 16841, 16841, 16841, 16817, 16817, 16817, 16788, 16788, 16788, 16764, 16764, 16764, 16734, 16734, 16734, 16710, 16710, 16680, 16680, 16680, 16657, 16657, 16657, 16627, 16627, 16627, 16603, 16603, 16603, 16573, 16573, 16573, 16549, 16549, 16549, 16519, 16519, 16519, 16495, 16495, 16495, 16465, 16465, 16465, 16442, 16442, 16442, 16412, 16412, 16388, 16388, 16388, 16358, 16358, 16358, 16334, 16334, 16334, 16304, 16304, 16304, 16280, 16280, 16280, 16250, 16250, 16250, 16226, 16226, 16226, 16196, 16196, 16196, 16172, 16172, 16172, 16142, 16142, 16142, 16118, 16118, 16118, 16088, 16088, 16064, 16064, 16064, 16034, 16034, 16034, 16010, 16010, 16010, 15980, 15980, 15980, 15956, 15956, 15956, 15926, 15926, 15926, 15902, 15902, 15902, 15872, 15872, 15872, 15848, 15848, 15848, 15818, 15818, 15818, 15794, 15794, 15794, 15764, 15764, 15740, 15740, 15740, 15716, 15716, 15716, 15686, 15686, 15686, 15662, 15662, 15662, 15632, 15632, 15632, 15608, 15608, 15608, 15577, 15577, 15577, 15553, 15553, 15553, 15523, 15523, 15523, 15499, 15499, 15499, 15469, 15469, 15469, 15445, 15445, 15415, 15415, 15415, 15391, 15391, 15391, 15360, 15360, 15360, 15336, 15336, 15336, 15306, 15306, 15306, 15282, 15282, 15282, 15252, 15252, 15252, 15227, 15227, 15227, 15197, 15197, 15197, 15173, 15173, 15173, 15143, 15143, 15143, 15119, 15119, 15088, 15088, 15088, 15064, 15064, 15064, 15034, 15034, 15034, 15010, 15010, 15010, 14979, 14979, 14979, 14955, 14955, 14955, 14925, 14925, 14925, 14900, 14900, 14900, 14870, 14870, 14870, 14846, 14846, 14846, 14816, 14816, 14816, 14791, 14791, 14791, 14761, 14761, 14737, 14737, 14737, 14706, 14706, 14706, 14682, 14682, 14682, 14652, 14652, 14652, 14627, 14627, 14627, 14597, 14597, 14597, 14572, 14572, 14572, 14542, 14542, 14542, 14518, 14518, 14518, 14493, 14493, 14493, 14463, 14463, 14463, 14439, 14439, 14439, 14408, 14408, 14384, 14384, 14384, 14353, 14353, 14353, 14329, 14329, 14329, 14298, 14298, 14298, 14274, 14274, 14274, 14243, 14243, 14243, 14219, 14219, 14219, 14188, 14188, 14188, 14164, 14164, 14164, 14133, 14133, 14133, 14109, 14109, 14109, 14078, 14078, 14078, 14054, 14054, 14023, 14023, 14023, 13999, 13999, 13999, 13968, 13968, 13968, 13944, 13944, 13944, 13913, 13913, 13913, 13889, 13889, 13889, 13858, 13858, 13858, 13834, 13834, 13834, 13803, 13803, 13803, 13778, 13778, 13778, 13748, 13748, 13748, 13723, 13723, 13723, 13693, 13693, 13693, 13668, 13668, 13637, 13637, 13637, 13613, 13613, 13613, 13582, 13582, 13582, 13557, 13557, 13557, 13527, 13527, 13527, 13502, 13502, 13502, 13471, 13471, 13471, 13447, 13447, 13447, 13416, 13416, 13416, 13391, 13391, 13391, 13361, 13361, 13361, 13336, 13336, 13336, 13305, 13305, 13305, 13280, 13280, 13256, 13256, 13256, 13225, 13225, 13225, 13200, 13200, 13200, 13169, 13169, 13169, 13145, 13145, 13145, 13114, 13114, 13114, 13089, 13089, 13089, 13058, 13058, 13058, 13034, 13034, 13034, 13003, 13003, 13003, 12978, 12978, 12978, 12947, 12947, 12947, 12922, 12922, 12922, 12891, 12891, 12891, 12867, 12867, 12836, 12836, 12836, 12811, 12811, 12811, 12780, 12780, 12780, 12755, 12755, 12755, 12724, 12724, 12724, 12699, 12699, 12699, 12668, 12668, 12668, 12643, 12643, 12643, 12612, 12612, 12612, 12588, 12588, 12588, 12557, 12557, 12557, 12532, 12532, 12532, 12501, 12501, 12501, 12476, 12476, 12476, 12445, 12445, 12445, 12420, 12420, 12389, 12389, 12389, 12364, 12364, 12364, 12333, 12333, 12333, 12308, 12308, 12308, 12277, 12277, 12277, 12252, 12252, 12252, 12221, 12221, 12221, 12196, 12196, 12196, 12164, 12164, 12164, 12139, 12139, 12139, 12108, 12108, 12108, 12083, 12083, 12083, 12058, 12058, 12058, 12027, 12027, 12027, 12002, 12002, 12002, 11971, 11971, 11946, 11946, 11946, 11915, 11915, 11915, 11890, 11890, 11890, 11858, 11858, 11858, 11833, 11833, 11833, 11802, 11802, 11802, 11777, 11777, 11777, 11746, 11746, 11746, 11721, 11721, 11721, 11689, 11689, 11689, 11664, 11664, 11664, 11633, 11633, 11633, 11608, 11608, 11608, 11576, 11576, 11576, 11551, 11551, 11551, 11520, 11520, 11520, 11495, 11495, 11463, 11463, 11463, 11438, 11438, 11438, 11407, 11407, 11407, 11382, 11382, 11382, 11350, 11350, 11350, 11325, 11325, 11325, 11293, 11293, 11293, 11268, 11268, 11268, 11237, 11237, 11237, 11212, 11212, 11212, 11180, 11180, 11180, 11155, 11155, 11155, 11123, 11123, 11123, 11098, 11098, 11098, 11067, 11067, 11067, 11041, 11041, 11041, 11010, 11010, 10984, 10984, 10984, 10953, 10953, 10953, 10928, 10928, 10928, 10896, 10896, 10896, 10871, 10871, 10871, 10839, 10839, 10839, 10814, 10814, 10814, 10788, 10788, 10788, 10757, 10757, 10757, 10731, 10731, 10731, 10700, 10700, 10700, 10674, 10674, 10674, 10643, 10643, 10643, 10617, 10617, 10617, 10586, 10586, 10586, 10560, 10560, 10560, 10528, 10528, 10528, 10503, 10503, 10503, 10471, 10471, 10446, 10446, 10446, 10414, 10414, 10414, 10389, 10389, 10389, 10357, 10357, 10357, 10331, 10331, 10331, 10300, 10300, 10300, 10274, 10274, 10274, 10242, 10242, 10242, 10217, 10217, 10217, 10185, 10185, 10185, 10159, 10159, 10159, 10128, 10128, 10128, 10102, 10102, 10102, 10070, 10070, 10070, 10045, 10045, 10045, 10013, 10013, 10013, 9987, 9987, 9987, 9955, 9955, 9955, 9930, 9930, 9930, 9898, 9898, 9898, 9872, 9872, 9840, 9840, 9840, 9814, 9814, 9814, 9782, 9782, 9782, 9757, 9757, 9757, 9725, 9725, 9725, 9699, 9699, 9699, 9667, 9667, 9667, 9641, 9641, 9641, 9609, 9609, 9609, 9584, 9584, 9584, 9552, 9552, 9552, 9526, 9526, 9526, 9500, 9500, 9500, 9468, 9468, 9468, 9442, 9442, 9442, 9410, 9410, 9410, 9385, 9385, 9385, 9352, 9352, 9352, 9327, 9327, 9327, 9294, 9294, 9294, 9269, 9269, 9269, 9236, 9236, 9236, 9211, 9211, 9178, 9178, 9178, 9153, 9153, 9153, 9120, 9120, 9120, 9095, 9095, 9095, 9062, 9062, 9062, 9036, 9036, 9036, 9004, 9004, 9004, 8978, 8978, 8978, 8946, 8946, 8946, 8920, 8920, 8920, 8888, 8888, 8888, 8862, 8862, 8862, 8830, 8830, 8830, 8804, 8804, 8804, 8771, 8771, 8771, 8745, 8745, 8745, 8713, 8713, 8713, 8687, 8687, 8687, 8655, 8655, 8655, 8629, 8629, 8629, 8596, 8596, 8596, 8570, 8570, 8570, 8538, 8538, 8538, 8512, 8512, 8512, 8479, 8479, 8453, 8453, 8453, 8421, 8421, 8421, 8395, 8395, 8395, 8362, 8362, 8362, 8336, 8336, 8336, 8303, 8303, 8303, 8277, 8277, 8277, 8245, 8245, 8245, 8219, 8219, 8219, 8193, 8193, 8193, 8160, 8160, 8160, 8134, 8134, 8134, 8101, 8101, 8101, 8075, 8075, 8075, 8042, 8042, 8042, 8016, 8016, 8016, 7984, 7984, 7984, 7957, 7957, 7957, 7925, 7925, 7925, 7899, 7899, 7899, 7866, 7866, 7866, 7840, 7840, 7840, 7807, 7807, 7807, 7781, 7781, 7781, 7748, 7748, 7748, 7722, 7722, 7722, 7689, 7689, 7689, 7663, 7663, 7663, 7630, 7630, 7630, 7603, 7603, 7571, 7571, 7571, 7544, 7544, 7544, 7511, 7511, 7511, 7485, 7485, 7485, 7452, 7452, 7452, 7426, 7426, 7426, 7393, 7393, 7393, 7367, 7367, 7367, 7334, 7334, 7334, 7307, 7307, 7307, 7274, 7274, 7274, 7248, 7248, 7248, 7215, 7215, 7215, 7188, 7188, 7188, 7155, 7155, 7155, 7129, 7129, 7129, 7096, 7096, 7096, 7070, 7070, 7070, 7036, 7036, 7036, 7010, 7010, 7010, 6977, 6977, 6977, 6950, 6950, 6950, 6924, 6924, 6924, 6891, 6891, 6891, 6864, 6864, 6864, 6831, 6831, 6831, 6805, 6805, 6805, 6771, 6771, 6771, 6745, 6745, 6745, 6712, 6712, 6712, 6685, 6685, 6685, 6652, 6652, 6652, 6625, 6625, 6625, 6592, 6592, 6592, 6565, 6565, 6565, 6532, 6532, 6532, 6506, 6506, 6506, 6472, 6472, 6446, 6446, 6446, 6412, 6412, 6412, 6386, 6386, 6386, 6352, 6352, 6352, 6326, 6326, 6326, 6292, 6292, 6292, 6265, 6265, 6265, 6232, 6232, 6232, 6205, 6205, 6205, 6172, 6172, 6172, 6145, 6145, 6145, 6112, 6112, 6112, 6085, 6085, 6085, 6051, 6051, 6051, 6025, 6025, 6025, 5991, 5991, 5991, 5964, 5964, 5964, 5931, 5931, 5931, 5904, 5904, 5904, 5870, 5870, 5870, 5844, 5844, 5844, 5810, 5810, 5810, 5783, 5783, 5783, 5750, 5750, 5750, 5723, 5723, 5723, 5689, 5689, 5689, 5662, 5662, 5662, 5628, 5628, 5628, 5601, 5601, 5601, 5575, 5575, 5575, 5541, 5541, 5541, 5514, 5514, 5514, 5480, 5480, 5480, 5453, 5453, 5453, 5419, 5419, 5419, 5392, 5392, 5392, 5359, 5359, 5359, 5332, 5332, 5332, 5298, 5298, 5298, 5271, 5271, 5271, 5237, 5237, 5237, 5210, 5210, 5210, 5176, 5176, 5176, 5149, 5149, 5149, 5115, 5115, 5115, 5088, 5088, 5088, 5054, 5054, 5054, 5027, 5027, 5027, 4993, 4993, 4993, 4966, 4966, 4966, 4932, 4932, 4932, 4905, 4905, 4905, 4871, 4871, 4871, 4844, 4844, 4844, 4810, 4810, 4810, 4782, 4782, 4782, 4748, 4748, 4748, 4721, 4721, 4721, 4687, 4687, 4687, 4660, 4660, 4660, 4626, 4626, 4626, 4598, 4598, 4598, 4564, 4564, 4564, 4537, 4537, 4537, 4503, 4503, 4503, 4475, 4475, 4475, 4441, 4441, 4441, 4414, 4414, 4414, 4380, 4380, 4380, 4352, 4352, 4352, 4318, 4318, 4318, 4291, 4291, 4291, 4257, 4257, 4257, 4229, 4229, 4229, 4202, 4202, 4202, 4167, 4167, 4167, 4140, 4140, 4140, 4106, 4106, 4106, 4078, 4078, 4078, 4044, 4044, 4016, 4016, 4016, 3982, 3982, 3982, 3954, 3954, 3954, 3920, 3920, 3920, 3893, 3893, 3893, 3858, 3858, 3858, 3831, 3831, 3831, 3796, 3796, 3796, 3769, 3769, 3769, 3734, 3734, 3734, 3706, 3706, 3706, 3672, 3672, 3672, 3644, 3644, 3644, 3610, 3610, 3610, 3582, 3582, 3582, 3548, 3548, 3548, 3520, 3520, 3520, 3485, 3485, 3485, 3458, 3458, 3458, 3423, 3423, 3423, 3395, 3395, 3395, 3361, 3361, 3361, 3333, 3333, 3333, 3298, 3298, 3298, 3298, 3270, 3270, 3270, 3236, 3236, 3236, 3208, 3208, 3208, 3173, 3173, 3173, 3145, 3145, 3145, 3111, 3111, 3111, 3083, 3083, 3083, 3048, 3048, 3048, 3020, 3020, 3020, 2985, 2985, 2985, 2957, 2957, 2957, 2923, 2923, 2923, 2895, 2895, 2895, 2860, 2860, 2860, 2832, 2832, 2832, 2804, 2804, 2804, 2769, 2769, 2769, 2741, 2741, 2741, 2706, 2706, 2706, 2678, 2678, 2678, 2643, 2643, 2643, 2615, 2615, 2615, 2580, 2580, 2580, 2552, 2552, 2552, 2517, 2517, 2517, 2489, 2489, 2489, 2454, 2454, 2454, 2426, 2426, 2426, 2391, 2391, 2391, 2363, 2363, 2363, 2328, 2328, 2328, 2299, 2299, 2299, 2264, 2264, 2264, 2236, 2236, 2236, 2201, 2201, 2201, 2173, 2173, 2173, 2138, 2138, 2138, 2109, 2109, 2109, 2074, 2074, 2074, 2046, 2046, 2046, 2011, 2011, 2011, 1982, 1982, 1982, 1947, 1947, 1947, 1919, 1919, 1919, 1883, 1883, 1883, 1855, 1855, 1855, 1820, 1820, 1820, 1792, 1792, 1792, 1756, 1756, 1756, 1728, 1728, 1728, 1692, 1692, 1692, 1664, 1664, 1664, 1629, 1629, 1629, 1600, 1600, 1600, 1565, 1565, 1565, 1536, 1536, 1536, 1501, 1501, 1501, 1472, 1472, 1472, 1437, 1437, 1437, 1408, 1408, 1408, 1380, 1380, 1380, 1344, 1344, 1344, 1316, 1316, 1316, 1280, 1280, 1280, 1252, 1252, 1252, 1216, 1216, 1216, 1187, 1187, 1187, 1152, 1152, 1152, 1123, 1123, 1123, 1087, 1087, 1087, 1059, 1059, 1059, 1023, 1023, 1023, 994, 994, 994, 959, 959, 959, 930, 930, 930, 894, 894, 894, 894, 865, 865, 865, 830, 830, 830, 801, 801, 801, 765, 765, 765, 736, 736, 736, 700, 700, 700, 672, 672, 672, 636, 636, 636, 607, 607, 607, 571, 571, 571, 542, 542, 542, 506, 506, 506, 477, 477, 477, 441, 441, 441, 412, 412, 412, 376, 376, 376, 347, 347, 347, 311, 311, 311, 282, 282, 282, 246, 246, 246, 217, 217, 217, 181, 181, 181, 152, 152, 152, 116, 116, 116, 87, 87, 87, 51, 51, 51, 22, 22, 22, 71993, 71993, 71993, 71956, 71956, 71956, 71927, 71927, 71927, 71891, 71891, 71891, 71862, 71862, 71862, 71826, 71826, 71826, 71797, 71797, 71797, 71761, 71761, 71761, 71732, 71732, 71732, 71732, 71696, 71696, 71696, 71667, 71667, 71667, 71631, 71631, 71631, 71602, 71602, 71602, 71566, 71566, 71566, 71537, 71537, 71537, 71501, 71501, 71501, 71472, 71472, 71472, 71436, 71436, 71436, 71408, 71408, 71408, 71372, 71372, 71372, 71343, 71343, 71343, 71307, 71307, 71307, 71278, 71278, 71278, 71242, 71242, 71242, 71213, 71213, 71213, 71178, 71178, 71178, 71149, 71149, 71149, 71113, 71113, 71113, 71084, 71084, 71084, 71049, 71049, 71049, 71020, 71020, 71020, 70984, 70984, 70984, 70956, 70956, 70956, 70920, 70920, 70920, 70891, 70891, 70891, 70856, 70856, 70856, 70856, 70827, 70827, 70827, 70791, 70791, 70791, 70763, 70763, 70763, 70727, 70727, 70727, 70699, 70699, 70699, 70663, 70663, 70663, 70634, 70634, 70634, 70599, 70599, 70599, 70570, 70570, 70570, 70542, 70542, 70542, 70506, 70506, 70506, 70478, 70478, 70478, 70442, 70442, 70442, 70414, 70414, 70414, 70379, 70379, 70379, 70350, 70350, 70350, 70315, 70315, 70315, 70286, 70286, 70286, 70251, 70251, 70251, 70223, 70223, 70223, 70187, 70187, 70187, 70159, 70159, 70159, 70159, 70124, 70124, 70124, 70095, 70095, 70095, 70060, 70060, 70060, 70032, 70032, 70032, 69996, 69996, 69996, 69968, 69968, 69968, 69933, 69933, 69933, 69905, 69905, 69905, 69869, 69869, 69869, 69841, 69841, 69841, 69806, 69806, 69806, 69778, 69778, 69778, 69743, 69743, 69743, 69715, 69715, 69715, 69679, 69679, 69679, 69651, 69651, 69651, 69616, 69616, 69616, 69588, 69588, 69588, 69553, 69553, 69553, 69525, 69525, 69525, 69525, 69490, 69490, 69490, 69462, 69462, 69462, 69427, 69427, 69427, 69399, 69399, 69399, 69364, 69364, 69364, 69336, 69336, 69336, 69301, 69301, 69301, 69273, 69273, 69273, 69238, 69238, 69238, 69210, 69210, 69210, 69175, 69175, 69175, 69147, 69147, 69147, 69119, 69119, 69119, 69084, 69084, 69084, 69056, 69056, 69056, 69022, 69022, 69022, 68994, 68994, 68994, 68959, 68959, 68959, 68959, 68931, 68931, 68931, 68896, 68896, 68896, 68868, 68868, 68868, 68834, 68834, 68834, 68806, 68806, 68806, 68771, 68771, 68771, 68743, 68743, 68743, 68709, 68709, 68709, 68681, 68681, 68681, 68646, 68646, 68646, 68619, 68619, 68619, 68584, 68584, 68584, 68556, 68556, 68556, 68522, 68522, 68522, 68494, 68494, 68494, 68459, 68459, 68459, 68459, 68432, 68432, 68432, 68397, 68397, 68397, 68369, 68369, 68369, 68335, 68335, 68335, 68307, 68307, 68307, 68273, 68273, 68273, 68245, 68245, 68245, 68211, 68211, 68211, 68183, 68183, 68183, 68149, 68149, 68149, 68121, 68121, 68121, 68087, 68087, 68087, 68059, 68059, 68059, 68025, 68025, 68025, 67997, 67997, 67997, 67997, 67963, 67963, 67963, 67936, 67936, 67936, 67901, 67901, 67901, 67874, 67874, 67874, 67839, 67839, 67839, 67812, 67812, 67812, 67778, 67778, 67778, 67750, 67750, 67750, 67723, 67723, 67723, 67689, 67689, 67689, 67661, 67661, 67661, 67627, 67627, 67627, 67600, 67600, 67600, 67566, 67566, 67566, 67566, 67538, 67538, 67538, 67504, 67504, 67504, 67477, 67477, 67477, 67443, 67443, 67443, 67415, 67415, 67415, 67381, 67381, 67381, 67354, 67354, 67354, 67320, 67320, 67320, 67293, 67293, 67293, 67259, 67259, 67259, 67231, 67231, 67231, 67197, 67197, 67197, 67170, 67170, 67170, 67170, 67136, 67136, 67136, 67109, 67109, 67109, 67075, 67075, 67075, 67048, 67048, 67048, 67014, 67014, 67014, 66987, 66987, 66987, 66953, 66953, 66953, 66926, 66926, 66926, 66892, 66892, 66892, 66865, 66865, 66865, 66831, 66831, 66831, 66804, 66804, 66804, 66804, 66770, 66770, 66770, 66743, 66743, 66743, 66709, 66709, 66709, 66682, 66682, 66682, 66648, 66648, 66648, 66621, 66621, 66621, 66587, 66587, 66587, 66560, 66560, 66560, 66527, 66527, 66527, 66500, 66500, 66500, 66466, 66466, 66466, 66439, 66439, 66439, 66439, 66412, 66412, 66412, 66378, 66378, 66378, 66351, 66351, 66351, 66318, 66318, 66318, 66291, 66291, 66291, 66257, 66257, 66257, 66230, 66230, 66230, 66197, 66197, 66197, 66170, 66170, 66170, 66136, 66136, 66136, 66109, 66109, 66109, 66076, 66076, 66076, 66076, 66049, 66049, 66049, 66016, 66016, 66016, 65989, 65989, 65989, 65955, 65955, 65955, 65928, 65928, 65928, 65895, 65895, 65895, 65868, 65868, 65868, 65835, 65835, 65835, 65808, 65808, 65808, 65775, 65775, 65775, 65748, 65748, 65748, 65748, 65715, 65715, 65715, 65688, 65688, 65688, 65654, 65654, 65654, 65628, 65628, 65628, 65594, 65594, 65594, 65568, 65568, 65568, 65534, 65534, 65534, 65508, 65508, 65508, 65475, 65475, 65475, 65448, 65448, 65448, 65448, 65415, 65415, 65415, 65388, 65388, 65388, 65355, 65355, 65355, 65328, 65328, 65328, 65295, 65295, 65295, 65268, 65268, 65268, 65235, 65235, 65235, 65209, 65209, 65209, 65175, 65175, 65175, 65149, 65149, 65149, 65149, 65116, 65116, 65116, 65089, 65089, 65089, 65063, 65063, 65063, 65030, 65030, 65030, 65003, 65003, 65003, 64970, 64970, 64970, 64944, 64944, 64944, 64911, 64911, 64911, 64884, 64884, 64884, 64851, 64851, 64851, 64851, 64825, 64825, 64825, 64792, 64792, 64792, 64765, 64765, 64765, 64732, 64732, 64732, 64706, 64706, 64706, 64673, 64673, 64673, 64647, 64647, 64647, 64614, 64614, 64614, 64587, 64587, 64587, 64587, 64554, 64554, 64554, 64528, 64528, 64528, 64495, 64495, 64495, 64469, 64469, 64469, 64436, 64436, 64436, 64410, 64410, 64410, 64377, 64377, 64377, 64351, 64351, 64351, 64318, 64318, 64318, 64318, 64292, 64292, 64292, 64259, 64259, 64259, 64232, 64232, 64232, 64200, 64200, 64200, 64173, 64173, 64173, 64141, 64141, 64141, 64115, 64115, 64115, 64082, 64082, 64082, 64056, 64056, 64056, 64056, 64023, 64023, 64023, 63997, 63997, 63997, 63964, 63964, 63964, 63938, 63938, 63938, 63905, 63905, 63905, 63879, 63879, 63879, 63847, 63847, 63847, 63820, 63820, 63820, 63788, 63788, 63788, 63788, 63762, 63762, 63762, 63736, 63736, 63736, 63703, 63703, 63703, 63677, 63677, 63677, 63644, 63644, 63644, 63618, 63618, 63618, 63586, 63586, 63586, 63560, 63560, 63560, 63560, 63527, 63527, 63527, 63501, 63501, 63501, 63469, 63469, 63469, 63443, 63443, 63443, 63410, 63410, 63410, 63384, 63384, 63384, 63352, 63352, 63352, 63326, 63326, 63326, 63326, 63294, 63294, 63294, 63268, 63268, 63268, 63235, 63235, 63235, 63209, 63209, 63209, 63177, 63177, 63177, 63151, 63151, 63151, 63119, 63119, 63119, 63093, 63093, 63093, 63093, 63060, 63060, 63060, 63035, 63035, 63035, 63002, 63002, 63002, 62976, 62976, 62976, 62944, 62944, 62944, 62918, 62918, 62918, 62886, 62886, 62886, 62860, 62860, 62860, 62860, 62828, 62828, 62828, 62802, 62802, 62802, 62770, 62770, 62770, 62744, 62744, 62744, 62712, 62712, 62712, 62686, 62686, 62686, 62654, 62654, 62654, 62628, 62628, 62628, 62628, 62596, 62596, 62596, 62570, 62570, 62570, 62538, 62538, 62538, 62513, 62513, 62513, 62480, 62480, 62480, 62455, 62455, 62455, 62429, 62429, 62429, 62429, 62397, 62397, 62397, 62371, 62371, 62371, 62339, 62339, 62339, 62314, 62314, 62314, 62282, 62282, 62282, 62256, 62256, 62256, 62224, 62224, 62224, 62198, 62198, 62198, 62198, 62166, 62166, 62166, 62141, 62141, 62141, 62109, 62109, 62109, 62083, 62083, 62083, 62051, 62051, 62051, 62026, 62026, 62026, 61994, 61994, 61994, 61994, 61968, 61968, 61968, 61936, 61936, 61936, 61911, 61911, 61911, 61879, 61879, 61879, 61853, 61853, 61853, 61821, 61821, 61821, 61796, 61796, 61796, 61796, 61764, 61764, 61764, 61739, 61739, 61739, 61707, 61707, 61707, 61681, 61681, 61681, 61649, 61649, 61649, 61624, 61624, 61624, 61592, 61592, 61592, 61592, 61567, 61567, 61567, 61535, 61535, 61535, 61510, 61510, 61510, 61478, 61478, 61478, 61452, 61452, 61452, 61421, 61421, 61421, 61421, 61395, 61395, 61395, 61364, 61364, 61364, 61338, 61338, 61338, 61307, 61307, 61307, 61281, 61281, 61281, 61250, 61250, 61250, 61224, 61224, 61224, 61224, 61193, 61193, 61193, 61167, 61167, 61167, 61142, 61142, 61142, 61110, 61110, 61110, 61085, 61085, 61085, 61053, 61053, 61053, 61028, 61028, 61028, 61028, 60997, 60997, 60997, 60971, 60971, 60971, 60940, 60940, 60940, 60915, 60915, 60915, 60883, 60883, 60883, 60858, 60858, 60858, 60858, 60826, 60826, 60826, 60801, 60801, 60801, 60769, 60769, 60769, 60744, 60744, 60744, 60713, 60713, 60713, 60688, 60688, 60688, 60688, 60656, 60656, 60656, 60631, 60631, 60631, 60600, 60600, 60600, 60574, 60574, 60574, 60543, 60543, 60543, 60518, 60518, 60518, 60486, 60486, 60486, 60486, 60461, 60461, 60461, 60430, 60430, 60430, 60405, 60405, 60405, 60373, 60373, 60373, 60348, 60348, 60348, 60317, 60317, 60317, 60317, 60292, 60292, 60292, 60261, 60261, 60261, 60236, 60236, 60236, 60204, 60204, 60204, 60179, 60179, 60179, 60148, 60148, 60148, 60148, 60123, 60123, 60123, 60092, 60092, 60092, 60067, 60067, 60067, 60035, 60035, 60035, 60010, 60010, 60010, 59979, 59979, 59979, 59979, 59954, 59954, 59954, 59929, 59929, 59929, 59898, 59898, 59898, 59873, 59873, 59873, 59842, 59842, 59842, 59842, 59817, 59817, 59817, 59786, 59786, 59786, 59761, 59761, 59761, 59730, 59730, 59730, 59705, 59705, 59705, 59674, 59674, 59674, 59674, 59649, 59649, 59649, 59618, 59618, 59618, 59593, 59593, 59593, 59562, 59562, 59562, 59537, 59537, 59537, 59506, 59506, 59506, 59506, 59481, 59481, 59481, 59450, 59450, 59450, 59425, 59425, 59425, 59394, 59394, 59394, 59369, 59369, 59369, 59369, 59338, 59338, 59338, 59313, 59313, 59313, 59282, 59282, 59282, 59257, 59257, 59257, 59226, 59226, 59226, 59202, 59202, 59202, 59202, 59171, 59171, 59171, 59146, 59146, 59146, 59115, 59115, 59115, 59090, 59090, 59090, 59059, 59059, 59059, 59059, 59034, 59034, 59034, 59004, 59004, 59004, 58979, 58979, 58979, 58948, 58948, 58948, 58923, 58923, 58923, 58892, 58892, 58892, 58892, 58868, 58868, 58868, 58837, 58837, 58837, 58812, 58812, 58812, 58781, 58781, 58781, 58757, 58757, 58757, 58757, 58726, 58726, 58726, 58701, 58701, 58701, 58676, 58676, 58676, 58646, 58646, 58646, 58621, 58621, 58621, 58621, 58590, 58590, 58590, 58566, 58566, 58566, 58535, 58535, 58535, 58510, 58510, 58510, 58479, 58479, 58479, 58455, 58455, 58455, 58455, 58424, 58424, 58424, 58400, 58400, 58400, 58369, 58369, 58369, 58344, 58344, 58344, 58314, 58314, 58314, 58314, 58289, 58289, 58289, 58258, 58258, 58258, 58234, 58234, 58234, 58203, 58203, 58203, 58179, 58179, 58179, 58179, 58148, 58148, 58148, 58124, 58124, 58124, 58093, 58093, 58093, 58068, 58068, 58068, 58038, 58038, 58038, 58038, 58013, 58013, 58013, 57983, 57983, 57983, 57958, 57958, 57958, 57928, 57928, 57928, 57903, 57903, 57903, 57903, 57873, 57873, 57873, 57848, 57848, 57848, 57818, 57818, 57818, 57793, 57793, 57793, 57763, 57763, 57763, 57763, 57738, 57738, 57738, 57708, 57708, 57708, 57683, 57683, 57683, 57653, 57653, 57653, 57629, 57629, 57629, 57629, 57598, 57598, 57598, 57574, 57574, 57574, 57543, 57543, 57543, 57519, 57519, 57519, 57519, 57488, 57488, 57488, 57464, 57464, 57464, 57440, 57440, 57440, 57409, 57409, 57409, 57385, 57385, 57385, 57385, 57355, 57355, 57355, 57330, 57330, 57330, 57300, 57300, 57300, 57276, 57276, 57276, 57245, 57245, 57245, 57245, 57221, 57221, 57221, 57191, 57191, 57191, 57166, 57166, 57166, 57136, 57136, 57136, 57136, 57112, 57112, 57112, 57081, 57081, 57081, 57057, 57057, 57057, 57027, 57027, 57027, 57003, 57003, 57003, 57003, 56972, 56972, 56972, 56948, 56948, 56948, 56918, 56918, 56918, 56894, 56894, 56894, 56863, 56863, 56863, 56863, 56839, 56839, 56839, 56809, 56809, 56809, 56785, 56785, 56785, 56754, 56754, 56754, 56754, 56730, 56730, 56730, 56700, 56700, 56700, 56676, 56676, 56676, 56646, 56646, 56646, 56622, 56622, 56622, 56622, 56591, 56591, 56591, 56567, 56567, 56567, 56537, 56537, 56537, 56513, 56513, 56513, 56513, 56483, 56483, 56483, 56459, 56459, 56459, 56429, 56429, 56429, 56404, 56404, 56404, 56404, 56374, 56374, 56374, 56350, 56350, 56350, 56320, 56320, 56320, 56296, 56296, 56296, 56266, 56266, 56266, 56266, 56242, 56242, 56242, 56218, 56218, 56218, 56188, 56188, 56188, 56164, 56164, 56164, 56164, 56134, 56134, 56134, 56110, 56110, 56110, 56080, 56080, 56080, 56056, 56056, 56056, 56056, 56026, 56026, 56026, 56002, 56002, 56002, 55972, 55972, 55972, 55948, 55948, 55948, 55918, 55918, 55918, 55918, 55894, 55894, 55894, 55864, 55864, 55864, 55840, 55840, 55840, 55810, 55810, 55810, 55810, 55786, 55786, 55786, 55756, 55756, 55756, 55732, 55732, 55732, 55702, 55702, 55702, 55702, 55678, 55678, 55678, 55648, 55648, 55648, 55624, 55624, 55624, 55594, 55594, 55594, 55594, 55570, 55570, 55570, 55541, 55541, 55541, 55517, 55517, 55517, 55487, 55487, 55487, 55487, 55463, 55463, 55463, 55433, 55433, 55433, 55409, 55409, 55409, 55379, 55379, 55379, 55379, 55355, 55355, 55355, 55326, 55326, 55326, 55302, 55302, 55302, 55272, 55272, 55272, 55272, 55248, 55248, 55248, 55218, 55218, 55218, 55194, 55194, 55194, 55165, 55165, 55165, 55165, 55141, 55141, 55141, 55111, 55111, 55111, 55087, 55087, 55087, 55063, 55063, 55063, 55063, 55034, 55034, 55034, 55010, 55010, 55010, 54980, 54980, 54980, 54956, 54956, 54956, 54956, 54927, 54927, 54927, 54903, 54903, 54903, 54873, 54873, 54873, 54849, 54849, 54849, 54849, 54820, 54820, 54820, 54796, 54796, 54796, 54766, 54766, 54766, 54743, 54743, 54743, 54743, 54713, 54713, 54713, 54689, 54689, 54689, 54660, 54660, 54660, 54636, 54636, 54636, 54636, 54606, 54606, 54606, 54583, 54583, 54583, 54553, 54553, 54553, 54529, 54529, 54529, 54529, 54500, 54500, 54500, 54476, 54476, 54476, 54446, 54446, 54446, 54446, 54423, 54423, 54423, 54393, 54393, 54393, 54369, 54369, 54369, 54340, 54340, 54340, 54340, 54316, 54316, 54316, 54287, 54287, 54287, 54263, 54263, 54263, 54234, 54234, 54234, 54234, 54210, 54210, 54210, 54180, 54180, 54180, 54157, 54157, 54157, 54127, 54127, 54127, 54127, 54104, 54104, 54104, 54074, 54074, 54074, 54051, 54051, 54051, 54051, 54021, 54021, 54021, 53998, 53998, 53998, 53968, 53968, 53968, 53944, 53944, 53944, 53944, 53915, 53915, 53915, 53891, 53891, 53891, 53868, 53868, 53868, 53838, 53838, 53838, 53838, 53815, 53815, 53815, 53785, 53785, 53785, 53762, 53762, 53762, 53762, 53733, 53733, 53733, 53709, 53709, 53709, 53680, 53680, 53680, 53656, 53656, 53656, 53656, 53627, 53627, 53627, 53603, 53603, 53603, 53574, 53574, 53574, 53574, 53550, 53550, 53550, 53521, 53521, 53521, 53498, 53498, 53498, 53468, 53468, 53468, 53468, 53445, 53445, 53445, 53415, 53415, 53415, 53392, 53392, 53392, 53392, 53363, 53363, 53363, 53339, 53339, 53339, 53310, 53310, 53310, 53286, 53286, 53286, 53286, 53257, 53257, 53257, 53234, 53234, 53234, 53204, 53204, 53204, 53204, 53181, 53181, 53181, 53152, 53152, 53152, 53128, 53128, 53128, 53099, 53099, 53099, 53099, 53076, 53076, 53076, 53046, 53046, 53046, 53023, 53023, 53023, 53023, 52994, 52994, 52994, 52970, 52970, 52970, 52941, 52941, 52941, 52918, 52918, 52918, 52918, 52889, 52889, 52889, 52865, 52865, 52865, 52836, 52836, 52836, 52836, 52813, 52813, 52813, 52783, 52783, 52783, 52760, 52760, 52760, 52760, 52731, 52731, 52731, 52708, 52708, 52708, 52684, 52684, 52684, 52655, 52655, 52655, 52655, 52632, 52632, 52632, 52603, 52603, 52603, 52579, 52579, 52579, 52579, 52550, 52550, 52550, 52527, 52527, 52527, 52498, 52498, 52498, 52498, 52475, 52475, 52475, 52445, 52445, 52445, 52422, 52422, 52422, 52393, 52393, 52393, 52393, 52370, 52370, 52370, 52341, 52341, 52341, 52318, 52318, 52318, 52318, 52288, 52288, 52288, 52265, 52265, 52265, 52236, 52236, 52236, 52236, 52213, 52213, 52213, 52184, 52184, 52184, 52161, 52161, 52161, 52161, 52132, 52132, 52132, 52108, 52108, 52108, 52079, 52079, 52079, 52079, 52056, 52056, 52056, 52027, 52027, 52027, 52004, 52004, 52004, 51975, 51975, 51975, 51975, 51952, 51952, 51952, 51923, 51923, 51923, 51900, 51900, 51900, 51900, 51871, 51871, 51871, 51847, 51847, 51847, 51818, 51818, 51818, 51818, 51795, 51795, 51795, 51766, 51766, 51766, 51743, 51743, 51743, 51743, 51714, 51714, 51714, 51691, 51691, 51691, 51662, 51662, 51662, 51662, 51639, 51639, 51639, 51610, 51610, 51610, 51587, 51587, 51587, 51587, 51558, 51558, 51558, 51535, 51535, 51535, 51512, 51512, 51512, 51512, 51483, 51483, 51483, 51460, 51460, 51460, 51431, 51431, 51431, 51431, 51408, 51408, 51408, 51379, 51379, 51379, 51356, 51356, 51356, 51356, 51327, 51327, 51327, 51304, 51304, 51304, 51275, 51275, 51275, 51252, 51252, 51252, 51252, 51223, 51223, 51223, 51200, 51200, 51200, 51171, 51171, 51171, 51171, 51148, 51148, 51148, 51120, 51120, 51120, 51096, 51096, 51096, 51096, 51068, 51068, 51068, 51045, 51045, 51045, 51016, 51016, 51016, 51016, 50993, 50993, 50993, 50964, 50964, 50964, 50964, 50941, 50941, 50941, 50912, 50912, 50912, 50889, 50889, 50889, 50889, 50861, 50861, 50861, 50838, 50838, 50838, 50809, 50809, 50809, 50809, 50786, 50786, 50786, 50757, 50757, 50757, 50734, 50734, 50734, 50734, 50705, 50705, 50705, 50682, 50682, 50682, 50654, 50654, 50654, 50654, 50631, 50631, 50631, 50602, 50602, 50602, 50579, 50579, 50579, 50579, 50550, 50550, 50550, 50527, 50527, 50527, 50499, 50499, 50499, 50499, 50476, 50476, 50476, 50447, 50447, 50447, 50424, 50424, 50424, 50424, 50396, 50396, 50396, 50373, 50373, 50373, 50350, 50350, 50350, 50350, 50321, 50321, 50321, 50298, 50298, 50298, 50269, 50269, 50269, 50269, 50247, 50247, 50247, 50218, 50218, 50218, 50218, 50195, 50195, 50195, 50166, 50166, 50166, 50144, 50144, 50144, 50144, 50115, 50115, 50115, 50092, 50092, 50092, 50063, 50063, 50063, 50063, 50041, 50041, 50041, 50012, 50012, 50012, 49989, 49989, 49989, 49989, 49961, 49961, 49961, 49938, 49938, 49938, 49938, 49909, 49909, 49909, 49886, 49886, 49886, 49858, 49858, 49858, 49858, 49835, 49835, 49835, 49806, 49806, 49806, 49784, 49784, 49784, 49784, 49755, 49755, 49755, 49732, 49732, 49732, 49704, 49704, 49704, 49704, 49681, 49681, 49681, 49652, 49652, 49652, 49652, 49630, 49630, 49630, 49601, 49601, 49601, 49578, 49578, 49578, 49578, 49550, 49550, 49550, 49527, 49527, 49527, 49498, 49498, 49498, 49498, 49476, 49476, 49476, 49447, 49447, 49447, 49424, 49424, 49424, 49424, 49396, 49396, 49396, 49373, 49373, 49373, 49373, 49345, 49345, 49345, 49322, 49322, 49322, 49294, 49294, 49294, 49294, 49271, 49271, 49271, 49248, 49248, 49248, 49248, 49220, 49220, 49220, 49197, 49197, 49197, 49168, 49168, 49168, 49168, 49146, 49146, 49146, 49117, 49117, 49117, 49095, 49095, 49095, 49095, 49066, 49066, 49066, 49043, 49043, 49043, 49043, 49015, 49015, 49015, 48992, 48992, 48992, 48964, 48964, 48964, 48964, 48941, 48941, 48941, 48913, 48913, 48913, 48890, 48890, 48890, 48890, 48862, 48862, 48862, 48839, 48839, 48839, 48839, 48811, 48811, 48811, 48788, 48788, 48788, 48760, 48760, 48760, 48760, 48737, 48737, 48737, 48709, 48709, 48709, 48709, 48686, 48686, 48686, 48658, 48658, 48658, 48635, 48635, 48635, 48635, 48607, 48607, 48607, 48584, 48584, 48584, 48584, 48556, 48556, 48556, 48533, 48533, 48533, 48505, 48505, 48505, 48505, 48482, 48482, 48482, 48454, 48454, 48454, 48454, 48431, 48431, 48431, 48403, 48403, 48403, 48380, 48380, 48380, 48380, 48352, 48352, 48352, 48329, 48329, 48329, 48329, 48301, 48301, 48301, 48279, 48279, 48279, 48250, 48250, 48250, 48250, 48228, 48228, 48228, 48199, 48199, 48199, 48199, 48177, 48177, 48177, 48149, 48149, 48149, 48126, 48126, 48126, 48126, 48103, 48103, 48103, 48075, 48075, 48075, 48075, 48053, 48053, 48053, 48024, 48024, 48024, 48002, 48002, 48002, 48002, 47974, 47974, 47974, 47951, 47951, 47951, 47951, 47923, 47923, 47923, 47900, 47900, 47900, 47872, 47872, 47872, 47872, 47850, 47850, 47850, 47821, 47821, 47821, 47821, 47799, 47799, 47799, 47771, 47771, 47771, 47771, 47748, 47748, 47748, 47720, 47720, 47720, 47697, 47697, 47697, 47697, 47669, 47669, 47669, 47647, 47647, 47647, 47647, 47619, 47619, 47619, 47596, 47596, 47596, 47568, 47568, 47568, 47568, 47545, 47545, 47545, 47517, 47517, 47517, 47517, 47495, 47495, 47495, 47467, 47467, 47467, 47467, 47444, 47444, 47444, 47416, 47416, 47416, 47393, 47393, 47393, 47393, 47365, 47365, 47365, 47343, 47343, 47343, 47343, 47315, 47315, 47315, 47292, 47292, 47292, 47292, 47264, 47264, 47264, 47242, 47242, 47242, 47214, 47214, 47214, 47214, 47191, 47191, 47191, 47163, 47163, 47163, 47163, 47141, 47141, 47141, 47113, 47113, 47113, 47113, 47090, 47090, 47090, 47062, 47062, 47062, 47040, 47040, 47040, 47040, 47011, 47011, 47011, 46989, 46989, 46989, 46989, 46967, 46967, 46967, 46939, 46939, 46939, 46939, 46916, 46916, 46916, 46888, 46888, 46888, 46888, 46866, 46866, 46866, 46838, 46838, 46838, 46815, 46815, 46815, 46815, 46787, 46787, 46787, 46765, 46765, 46765, 46765, 46737, 46737, 46737, 46714, 46714, 46714, 46714, 46686, 46686, 46686, 46664, 46664, 46664, 46664, 46636, 46636, 46636, 46614, 46614, 46614, 46586, 46586, 46586, 46586, 46563, 46563, 46563, 46535, 46535, 46535, 46535, 46513, 46513, 46513, 46485, 46485, 46485, 46485, 46462, 46462, 46462, 46434, 46434, 46434, 46434, 46412, 46412, 46412, 46384, 46384, 46384, 46362, 46362, 46362, 46362, 46334, 46334, 46334, 46311, 46311, 46311, 46311, 46283, 46283, 46283, 46261, 46261, 46261, 46261, 46233, 46233, 46233, 46211, 46211, 46211, 46211, 46183, 46183, 46183, 46161, 46161, 46161, 46161, 46133, 46133, 46133, 46110, 46110, 46110, 46110, 46082, 46082, 46082, 46060, 46060, 46060, 46032, 46032, 46032, 46032, 46010, 46010, 46010, 45982, 45982, 45982, 45982, 45960, 45960, 45960, 45932, 45932, 45932, 45932, 45909, 45909, 45909, 45881, 45881, 45881, 45881, 45859, 45859, 45859, 45837, 45837, 45837, 45837, 45809, 45809, 45809, 45787, 45787, 45787, 45787, 45759, 45759, 45759, 45736, 45736, 45736, 45736, 45709, 45709, 45709, 45686, 45686, 45686, 45658, 45658, 45658, 45658, 45636, 45636, 45636, 45608, 45608, 45608, 45608, 45586, 45586, 45586, 45558, 45558, 45558, 45558, 45536, 45536, 45536, 45508, 45508, 45508, 45508, 45486, 45486, 45486, 45458, 45458, 45458, 45458, 45436, 45436, 45436, 45408, 45408, 45408, 45408, 45386, 45386, 45386, 45358, 45358, 45358, 45358, 45336, 45336, 45336, 45308, 45308, 45308, 45308, 45285, 45285, 45285, 45258, 45258, 45258, 45258, 45235, 45235, 45235, 45208, 45208, 45208, 45208, 45185, 45185, 45185, 45158, 45158, 45158, 45158, 45135, 45135, 45135, 45108, 45108, 45108, 45108, 45085, 45085, 45085, 45058, 45058, 45058, 45058, 45035, 45035, 45035, 45008, 45008, 45008, 45008, 44985, 44985, 44985, 44958, 44958, 44958, 44958, 44935, 44935, 44935, 44908, 44908, 44908, 44908, 44885, 44885, 44885, 44858, 44858, 44858, 44858, 44835, 44835, 44835, 44808, 44808, 44808, 44808, 44785, 44785, 44785, 44763, 44763, 44763, 44763, 44736, 44736, 44736, 44713, 44713, 44713, 44713, 44686, 44686, 44686, 44663, 44663, 44663, 44663, 44636, 44636, 44636, 44613, 44613, 44613, 44613, 44586, 44586, 44586, 44564, 44564, 44564, 44564, 44536, 44536, 44536, 44514, 44514, 44514, 44514, 44486, 44486, 44486, 44464, 44464, 44464, 44464, 44436, 44436, 44436, 44414, 44414, 44414, 44414, 44386, 44386, 44386, 44364, 44364, 44364, 44364, 44336, 44336, 44336, 44314, 44314, 44314, 44314, 44287, 44287, 44287, 44264, 44264, 44264, 44264, 44237, 44237, 44237, 44215, 44215, 44215, 44215, 44187, 44187, 44187, 44165, 44165, 44165, 44165, 44137, 44137, 44137, 44115, 44115, 44115, 44115, 44087, 44087, 44087, 44065, 44065, 44065, 44065, 44037, 44037, 44037, 44015, 44015, 44015, 44015, 43988, 43988, 43988, 43966, 43966, 43966, 43966, 43938, 43938, 43938, 43916, 43916, 43916, 43916, 43888, 43888, 43888, 43888, 43866, 43866, 43866, 43838, 43838, 43838, 43838, 43816, 43816, 43816, 43789, 43789, 43789, 43789, 43767, 43767, 43767, 43739, 43739, 43739, 43739, 43717, 43717, 43717, 43689, 43689, 43689, 43689, 43667, 43667, 43667, 43645, 43645, 43645, 43645, 43617, 43617, 43617, 43595, 43595, 43595, 43595, 43568, 43568, 43568, 43546, 43546, 43546, 43546, 43518, 43518, 43518, 43518, 43496, 43496, 43496, 43468, 43468, 43468, 43468, 43446, 43446, 43446, 43419, 43419, 43419, 43419, 43397, 43397, 43397, 43369, 43369, 43369, 43369, 43347, 43347, 43347, 43319, 43319, 43319, 43319, 43297, 43297, 43297, 43270, 43270, 43270, 43270, 43248, 43248, 43248, 43248, 43220, 43220, 43220, 43198, 43198, 43198, 43198, 43170, 43170, 43170, 43148, 43148, 43148, 43148, 43121, 43121, 43121, 43099, 43099, 43099, 43099, 43071, 43071, 43071, 43049, 43049, 43049, 43049, 43022, 43022, 43022, 43022, 43000, 43000, 43000, 42972, 42972, 42972, 42972, 42950, 42950, 42950, 42922, 42922, 42922, 42922, 42900, 42900, 42900, 42873, 42873, 42873, 42873, 42851, 42851, 42851, 42823, 42823, 42823, 42823, 42801, 42801, 42801, 42801, 42774, 42774, 42774, 42752, 42752, 42752, 42752, 42724, 42724, 42724, 42702, 42702, 42702, 42702, 42675, 42675, 42675, 42653, 42653, 42653, 42653, 42625, 42625, 42625, 42625, 42603, 42603, 42603, 42576, 42576, 42576, 42576, 42554, 42554, 42554, 42532, 42532, 42532, 42532, 42504, 42504, 42504, 42482, 42482, 42482, 42482, 42455, 42455, 42455, 42455, 42433, 42433, 42433, 42405, 42405, 42405, 42405, 42383, 42383, 42383, 42356, 42356, 42356, 42356, 42334, 42334, 42334, 42306, 42306, 42306, 42306, 42284, 42284, 42284, 42284, 42257, 42257, 42257, 42235, 42235, 42235, 42235, 42207, 42207, 42207, 42185, 42185, 42185, 42185, 42158, 42158, 42158, 42158, 42136, 42136, 42136, 42108, 42108, 42108, 42108, 42086, 42086, 42086, 42059, 42059, 42059, 42059, 42037, 42037, 42037, 42009, 42009, 42009, 42009, 41988, 41988, 41988, 41988, 41960, 41960, 41960, 41938, 41938, 41938, 41938, 41911, 41911, 41911, 41889, 41889, 41889, 41889, 41861, 41861, 41861, 41861, 41839, 41839, 41839, 41812, 41812, 41812, 41812, 41790, 41790, 41790, 41762, 41762, 41762, 41762, 41740, 41740, 41740, 41740, 41713, 41713, 41713, 41691, 41691, 41691, 41691, 41664, 41664, 41664, 41642, 41642, 41642, 41642, 41614, 41614, 41614, 41614, 41592, 41592, 41592, 41565, 41565, 41565, 41565, 41543, 41543, 41543, 41516, 41516, 41516, 41516, 41494, 41494, 41494, 41494, 41466, 41466, 41466, 41444, 41444, 41444, 41444, 41422, 41422, 41422, 41395, 41395, 41395, 41395, 41373, 41373, 41373, 41373, 41346, 41346, 41346, 41324, 41324, 41324, 41324, 41296, 41296, 41296, 41296, 41274, 41274, 41274, 41247, 41247, 41247, 41247, 41225, 41225, 41225, 41198, 41198, 41198, 41198, 41176, 41176, 41176, 41176, 41148, 41148, 41148, 41126, 41126, 41126, 41126, 41099, 41099, 41099, 41099, 41077, 41077, 41077, 41050, 41050, 41050, 41050, 41028, 41028, 41028, 41000, 41000, 41000, 41000, 40979, 40979, 40979, 40979, 40951, 40951, 40951, 40929, 40929, 40929, 40929, 40902, 40902, 40902, 40902, 40880, 40880, 40880, 40853, 40853, 40853, 40853, 40831, 40831, 40831, 40803, 40803, 40803, 40803, 40781, 40781, 40781, 40781, 40754, 40754, 40754, 40732, 40732, 40732, 40732, 40705, 40705, 40705, 40705, 40683, 40683, 40683, 40656, 40656, 40656, 40656, 40634, 40634, 40634, 40634, 40606, 40606, 40606, 40584, 40584, 40584, 40584, 40557, 40557, 40557, 40535, 40535, 40535, 40535, 40508, 40508, 40508, 40508, 40486, 40486, 40486, 40459, 40459, 40459, 40459, 40437, 40437, 40437, 40437, 40409, 40409, 40409, 40388, 40388, 40388, 40388, 40360, 40360, 40360, 40360, 40338, 40338, 40338, 40316, 40316, 40316, 40316, 40289, 40289, 40289, 40289, 40267, 40267, 40267, 40240, 40240, 40240, 40240, 40218, 40218, 40218, 40218, 40191, 40191, 40191, 40169, 40169, 40169, 40169, 40142, 40142, 40142, 40142, 40120, 40120, 40120, 40092, 40092, 40092, 40092, 40070, 40070, 40070, 40070, 40043, 40043, 40043, 40021, 40021, 40021, 40021, 39994, 39994, 39994, 39994, 39972, 39972, 39972, 39945, 39945, 39945, 39945, 39923, 39923, 39923, 39923, 39896, 39896, 39896, 39874, 39874, 39874, 39874, 39846, 39846, 39846, 39846, 39825, 39825, 39825, 39797, 39797, 39797, 39797, 39775, 39775, 39775, 39775, 39748, 39748, 39748, 39726, 39726, 39726, 39726, 39699, 39699, 39699, 39699, 39677, 39677, 39677, 39650, 39650, 39650, 39650, 39628, 39628, 39628, 39628, 39601, 39601, 39601, 39579, 39579, 39579, 39579, 39552, 39552, 39552, 39552, 39530, 39530, 39530, 39502, 39502, 39502, 39502, 39481, 39481, 39481, 39481, 39453, 39453, 39453, 39432, 39432, 39432, 39432, 39404, 39404, 39404, 39404, 39382, 39382, 39382, 39355, 39355, 39355, 39355, 39333, 39333, 39333, 39333, 39306, 39306, 39306, 39284, 39284, 39284, 39284, 39262, 39262, 39262, 39262, 39235, 39235, 39235, 39235, 39213, 39213, 39213, 39186, 39186, 39186, 39186, 39164, 39164, 39164, 39164, 39137, 39137, 39137, 39115, 39115, 39115, 39115, 39088, 39088, 39088, 39088, 39066, 39066, 39066, 39039, 39039, 39039, 39039, 39017, 39017, 39017, 39017, 38990, 38990, 38990, 38990, 38968, 38968, 38968, 38941, 38941, 38941, 38941, 38919, 38919, 38919, 38919, 38891, 38891, 38891, 38870, 38870, 38870, 38870, 38842, 38842, 38842, 38842, 38821, 38821, 38821, 38821, 38793, 38793, 38793, 38771, 38771, 38771, 38771, 38744, 38744, 38744, 38744, 38722, 38722, 38722, 38695, 38695, 38695, 38695, 38673, 38673, 38673, 38673, 38646, 38646, 38646, 38646, 38624, 38624, 38624, 38597, 38597, 38597, 38597, 38575, 38575, 38575, 38575, 38548, 38548, 38548, 38526, 38526, 38526, 38526, 38499, 38499, 38499, 38499, 38477, 38477, 38477, 38477, 38450, 38450, 38450, 38428, 38428, 38428, 38428, 38401, 38401, 38401, 38401, 38379, 38379, 38379, 38352, 38352, 38352, 38352, 38330, 38330, 38330, 38330, 38303, 38303, 38303, 38303, 38281, 38281, 38281, 38254, 38254, 38254, 38254, 38232, 38232, 38232, 38232, 38205, 38205, 38205, 38205, 38183, 38183, 38183, 38161, 38161, 38161, 38161, 38134, 38134, 38134, 38134, 38112, 38112, 38112, 38112, 38085, 38085, 38085, 38063, 38063, 38063, 38063, 38036, 38036, 38036, 38036, 38014, 38014, 38014, 38014, 37987, 37987, 37987, 37965, 37965, 37965, 37965, 37938, 37938, 37938, 37938, 37916, 37916, 37916, 37916, 37889, 37889, 37889, 37867, 37867, 37867, 37867, 37840, 37840, 37840, 37840, 37818, 37818, 37818, 37818, 37791, 37791, 37791, 37769, 37769, 37769, 37769, 37742, 37742, 37742, 37742, 37720, 37720, 37720, 37720, 37693, 37693, 37693, 37671, 37671, 37671, 37671, 37644, 37644, 37644, 37644, 37622, 37622, 37622, 37622, 37595, 37595, 37595, 37573, 37573, 37573, 37573, 37546, 37546, 37546, 37546, 37524, 37524, 37524, 37524, 37497, 37497, 37497, 37475, 37475, 37475, 37475, 37448, 37448, 37448, 37448, 37426, 37426, 37426, 37426, 37399, 37399, 37399, 37377, 37377, 37377, 37377, 37350, 37350, 37350, 37350, 37328, 37328, 37328, 37328, 37301, 37301, 37301, 37301, 37279, 37279, 37279, 37252, 37252, 37252, 37252, 37230, 37230, 37230, 37230, 37203, 37203, 37203, 37203, 37181, 37181, 37181, 37154, 37154, 37154, 37154, 37132, 37132, 37132, 37132, 37105, 37105, 37105, 37105, 37083, 37083, 37083, 37083, 37061, 37061, 37061, 37034, 37034, 37034, 37034, 37012, 37012, 37012, 37012, 36985, 36985, 36985, 36985, 36963, 36963, 36963, 36963, 36936, 36936, 36936, 36914, 36914, 36914, 36914, 36887, 36887, 36887, 36887, 36865, 36865, 36865, 36865, 36838, 36838, 36838, 36816, 36816, 36816, 36816, 36789, 36789, 36789, 36789, 36767, 36767, 36767, 36767, 36740, 36740, 36740, 36740, 36718, 36718, 36718, 36691, 36691, 36691, 36691, 36669, 36669, 36669, 36669, 36642, 36642, 36642, 36642, 36620, 36620, 36620, 36620, 36593, 36593, 36593, 36593, 36571, 36571, 36571, 36544, 36544, 36544, 36544, 36522, 36522, 36522, 36522, 36495, 36495, 36495, 36495, 36473, 36473, 36473, 36473, 36446, 36446, 36446, 36424, 36424, 36424, 36424, 36397, 36397, 36397, 36397, 36375, 36375, 36375, 36375, 36348, 36348, 36348, 36348, 36326, 36326, 36326, 36299, 36299, 36299, 36299, 36278, 36278, 36278, 36278, 36250, 36250, 36250, 36250, 36229, 36229, 36229, 36229, 36201, 36201, 36201, 36201, 36180, 36180, 36180, 36152, 36152, 36152, 36152, 36131, 36131, 36131, 36131, 36103, 36103, 36103, 36103, 36082, 36082, 36082, 36082, 36054, 36054, 36054, 36054, 36033, 36033, 36033, 36005, 36005, 36005, 36005, 35984, 35984, 35984, 35984, 35962, 35962, 35962, 35962, 35935, 35935, 35935, 35935, 35913, 35913, 35913, 35913, 35886, 35886, 35886, 35864, 35864, 35864, 35864, 35837, 35837, 35837, 35837, 35815, 35815, 35815, 35815, 35788, 35788, 35788, 35788, 35766, 35766, 35766, 35766, 35739, 35739, 35739, 35717, 35717, 35717, 35717, 35690, 35690, 35690, 35690, 35668, 35668, 35668, 35668, 35641, 35641, 35641, 35641, 35619, 35619, 35619, 35619, 35592, 35592, 35592, 35592, 35570, 35570, 35570, 35543, 35543, 35543, 35543, 35521, 35521, 35521, 35521, 35494, 35494, 35494, 35494, 35472, 35472, 35472, 35472, 35445, 35445, 35445, 35445, 35423, 35423, 35423, 35423, 35396, 35396, 35396, 35374, 35374, 35374, 35374, 35347, 35347, 35347, 35347, 35325, 35325, 35325, 35325, 35298, 35298, 35298, 35298, 35276, 35276, 35276, 35276, 35249, 35249, 35249, 35249, 35227, 35227, 35227, 35200, 35200, 35200, 35200, 35178, 35178, 35178, 35178, 35151, 35151, 35151, 35151, 35129, 35129, 35129, 35129, 35102, 35102, 35102, 35102, 35080, 35080, 35080, 35080, 35053, 35053, 35053, 35053, 35031, 35031, 35031, 35031, 35004, 35004, 35004, 34982, 34982, 34982, 34982, 34955, 34955, 34955, 34955, 34933, 34933, 34933, 34933, 34912, 34912, 34912, 34912, 34884, 34884, 34884, 34884, 34863, 34863, 34863, 34863, 34835, 34835, 34835, 34835, 34814, 34814, 34814, 34786, 34786, 34786, 34786, 34765, 34765, 34765, 34765, 34737, 34737, 34737, 34737, 34716, 34716, 34716, 34716, 34688, 34688, 34688, 34688, 34667, 34667, 34667, 34667, 34639, 34639, 34639, 34639, 34618, 34618, 34618, 34618, 34590, 34590, 34590, 34590, 34569, 34569, 34569, 34541, 34541, 34541, 34541, 34520, 34520, 34520, 34520, 34492, 34492, 34492, 34492, 34471, 34471, 34471, 34471, 34443, 34443, 34443, 34443, 34422, 34422, 34422, 34422, 34394, 34394, 34394, 34394, 34373, 34373, 34373, 34373, 34345, 34345, 34345, 34345, 34324, 34324, 34324, 34324, 34296, 34296, 34296, 34275, 34275, 34275, 34275, 34247, 34247, 34247, 34247, 34226, 34226, 34226, 34226, 34198, 34198, 34198, 34198, 34177, 34177, 34177, 34177, 34149, 34149, 34149, 34149, 34128, 34128, 34128, 34128, 34100, 34100, 34100, 34100, 34079, 34079, 34079, 34079, 34051, 34051, 34051, 34051, 34030, 34030, 34030, 34030, 34002, 34002, 34002, 34002, 33981, 33981, 33981, 33981, 33953, 33953, 33953, 33932, 33932, 33932, 33932, 33904, 33904, 33904, 33904, 33882, 33882, 33882, 33882, 33855, 33855, 33855, 33855, 33833, 33833, 33833, 33833, 33812, 33812, 33812, 33812, 33784, 33784, 33784, 33784, 33763, 33763, 33763, 33763, 33735, 33735, 33735, 33735, 33714, 33714, 33714, 33714, 33686, 33686, 33686, 33686, 33665, 33665, 33665, 33665, 33637, 33637, 33637, 33637, 33616, 33616, 33616, 33616, 33588, 33588, 33588, 33588, 33566, 33566, 33566, 33566, 33539, 33539, 33539, 33539, 33517, 33517, 33517, 33517, 33490, 33490, 33490, 33468, 33468, 33468, 33468, 33441, 33441, 33441, 33441, 33419, 33419, 33419, 33419, 33392, 33392, 33392, 33392, 33370, 33370, 33370, 33370, 33343, 33343, 33343, 33343, 33321, 33321, 33321, 33321, 33294, 33294, 33294, 33294, 33272, 33272, 33272, 33272, 33245, 33245, 33245, 33245, 33223, 33223, 33223, 33223, 33196, 33196, 33196, 33196, 33174, 33174, 33174, 33174, 33147, 33147, 33147, 33147, 33125, 33125, 33125, 33125, 33098, 33098, 33098, 33098, 33076, 33076, 33076, 33076, 33049, 33049, 33049, 33049, 33027, 33027, 33027, 33027, 32999, 32999, 32999, 32999, 32978, 32978, 32978, 32978, 32950, 32950, 32950, 32950, 32929, 32929, 32929, 32929, 32901, 32901, 32901, 32901, 32879, 32879, 32879, 32879, 32852, 32852, 32852, 32852, 32830, 32830, 32830, 32830, 32803, 32803, 32803, 32803, 32781, 32781, 32781, 32781, 32754, 32754, 32754, 32754, 32732, 32732, 32732, 32732, 32710, 32710, 32710, 32710, 32683, 32683, 32683, 32683, 32661, 32661, 32661, 32661, 32634, 32634, 32634, 32634, 32612, 32612, 32612, 32612, 32585, 32585, 32585, 32585, 32563, 32563, 32563, 32563, 32536, 32536, 32536, 32536, 32514, 32514, 32514, 32514, 32487, 32487, 32487, 32487, 32465, 32465, 32465, 32465, 32437, 32437, 32437, 32437, 32416, 32416, 32416, 32416, 32388, 32388, 32388, 32388, 32366, 32366, 32366, 32366, 32339, 32339, 32339, 32339, 32317, 32317, 32317, 32317, 32290, 32290, 32290, 32290, 32268, 32268, 32268, 32268, 32241, 32241, 32241, 32241, 32219, 32219, 32219, 32219, 32192, 32192, 32192, 32192, 32170, 32170, 32170, 32170, 32143, 32143, 32143, 32143, 32121, 32121, 32121, 32121, 32093, 32093, 32093, 32093, 32072, 32072, 32072, 32072, 32044, 32044, 32044, 32044, 32044, 32022, 32022, 32022, 32022, 31995, 31995, 31995, 31995, 31973, 31973, 31973, 31973, 31946, 31946, 31946, 31946, 31924, 31924, 31924, 31924, 31897, 31897, 31897, 31897, 31875, 31875, 31875, 31875, 31848, 31848, 31848, 31848, 31826, 31826, 31826, 31826, 31798, 31798, 31798, 31798, 31776, 31776, 31776, 31776, 31749, 31749, 31749, 31749, 31727, 31727, 31727, 31727, 31700, 31700, 31700, 31700, 31678, 31678, 31678, 31678, 31651, 31651, 31651, 31651, 31629, 31629, 31629, 31629, 31607, 31607, 31607, 31607, 31580, 31580, 31580, 31580, 31580, 31558, 31558, 31558, 31558, 31530, 31530, 31530, 31530, 31509, 31509, 31509, 31509, 31481, 31481, 31481, 31481, 31459, 31459, 31459, 31459, 31432, 31432, 31432, 31432, 31410, 31410, 31410, 31410, 31383, 31383, 31383, 31383, 31361, 31361, 31361, 31361, 31333, 31333, 31333, 31333, 31312, 31312, 31312, 31312, 31284, 31284, 31284, 31284, 31262, 31262, 31262, 31262, 31262, 31235, 31235, 31235, 31235, 31213, 31213, 31213, 31213, 31186, 31186, 31186, 31186, 31164, 31164, 31164, 31164, 31136, 31136, 31136, 31136, 31115, 31115, 31115, 31115, 31087, 31087, 31087, 31087, 31065, 31065, 31065, 31065, 31038, 31038, 31038, 31038, 31016, 31016, 31016, 31016, 31016, 30989, 30989, 30989, 30989, 30967, 30967, 30967, 30967, 30939, 30939, 30939, 30939, 30917, 30917, 30917, 30917, 30890, 30890, 30890, 30890, 30868, 30868, 30868, 30868, 30841, 30841, 30841, 30841, 30819, 30819, 30819, 30819, 30791, 30791, 30791, 30791, 30791, 30769, 30769, 30769, 30769, 30742, 30742, 30742, 30742, 30720, 30720, 30720, 30720, 30693, 30693, 30693, 30693, 30671, 30671, 30671, 30671, 30643, 30643, 30643, 30643, 30622, 30622, 30622, 30622, 30594, 30594, 30594, 30594, 30572, 30572, 30572, 30572, 30572, 30545, 30545, 30545, 30545, 30523, 30523, 30523, 30523, 30501, 30501, 30501, 30501, 30473, 30473, 30473, 30473, 30452, 30452, 30452, 30452, 30424, 30424, 30424, 30424, 30402, 30402, 30402, 30402, 30402, 30375, 30375, 30375, 30375, 30353, 30353, 30353, 30353, 30325, 30325, 30325, 30325, 30303, 30303, 30303, 30303, 30276, 30276, 30276, 30276, 30254, 30254, 30254, 30254, 30227, 30227, 30227, 30227, 30227, 30205, 30205, 30205, 30205, 30177, 30177, 30177, 30177, 30155, 30155, 30155, 30155, 30128, 30128, 30128, 30128, 30106, 30106, 30106, 30106, 30078, 30078, 30078, 30078, 30078, 30056, 30056, 30056, 30056, 30029, 30029, 30029, 30029, 30007, 30007, 30007, 30007, 29980, 29980, 29980, 29980, 29958, 29958, 29958, 29958, 29930, 29930, 29930, 29930, 29930, 29908, 29908, 29908, 29908, 29881, 29881, 29881, 29881, 29859, 29859, 29859, 29859, 29831, 29831, 29831, 29831, 29809, 29809, 29809, 29809, 29782, 29782, 29782, 29782, 29782, 29760, 29760, 29760, 29760, 29732, 29732, 29732, 29732, 29710, 29710, 29710, 29710, 29683, 29683, 29683, 29683, 29661, 29661, 29661, 29661, 29661, 29633, 29633, 29633, 29633, 29611, 29611, 29611, 29611, 29584, 29584, 29584, 29584, 29562, 29562, 29562, 29562, 29534, 29534, 29534, 29534, 29534, 29512, 29512, 29512, 29512, 29485, 29485, 29485, 29485, 29463, 29463, 29463, 29463, 29441, 29441, 29441, 29441, 29413, 29413, 29413, 29413, 29413, 29391, 29391, 29391, 29391, 29364, 29364, 29364, 29364, 29342, 29342, 29342, 29342, 29314, 29314, 29314, 29314, 29292, 29292, 29292, 29292, 29292, 29265, 29265, 29265, 29265, 29243, 29243, 29243, 29243, 29215, 29215, 29215, 29215, 29193, 29193, 29193, 29193, 29166, 29166, 29166, 29166, 29166, 29144, 29144, 29144, 29144, 29116, 29116, 29116, 29116, 29094, 29094, 29094, 29094, 29066, 29066, 29066, 29066, 29066, 29044, 29044, 29044, 29044, 29017, 29017, 29017, 29017, 28995, 28995, 28995, 28995, 28967, 28967, 28967, 28967, 28967, 28945, 28945, 28945, 28945, 28918, 28918, 28918, 28918, 28896, 28896, 28896, 28896, 28868, 28868, 28868, 28868, 28846, 28846, 28846, 28846, 28846, 28818, 28818, 28818, 28818, 28796, 28796, 28796, 28796, 28769, 28769, 28769, 28769, 28747, 28747, 28747, 28747, 28747, 28719, 28719, 28719, 28719, 28697, 28697, 28697, 28697, 28670, 28670, 28670, 28670, 28648, 28648, 28648, 28648, 28648, 28620, 28620, 28620, 28620, 28598, 28598, 28598, 28598, 28570, 28570, 28570, 28570, 28570, 28548, 28548, 28548, 28548, 28521, 28521, 28521, 28521, 28499, 28499, 28499, 28499, 28471, 28471, 28471, 28471, 28471, 28449, 28449, 28449, 28449, 28421, 28421, 28421, 28421, 28399, 28399, 28399, 28399, 28372, 28372, 28372, 28372, 28372, 28349, 28349, 28349, 28349, 28327, 28327, 28327, 28327, 28300, 28300, 28300, 28300, 28300, 28278, 28278, 28278, 28278, 28250, 28250, 28250, 28250, 28228, 28228, 28228, 28228, 28200, 28200, 28200, 28200, 28200, 28178, 28178, 28178, 28178, 28151, 28151, 28151, 28151, 28128, 28128, 28128, 28128, 28128, 28101, 28101, 28101, 28101, 28079, 28079, 28079, 28079, 28051, 28051, 28051, 28051, 28029, 28029, 28029, 28029, 28029, 28001, 28001, 28001, 28001, 27979, 27979, 27979, 27979, 27951, 27951, 27951, 27951, 27951, 27929, 27929, 27929, 27929, 27902, 27902, 27902, 27902, 27880, 27880, 27880, 27880, 27880, 27852, 27852, 27852, 27852, 27830, 27830, 27830, 27830, 27802, 27802, 27802, 27802, 27802, 27780, 27780, 27780, 27780, 27752, 27752, 27752, 27752, 27730, 27730, 27730, 27730, 27730, 27702, 27702, 27702, 27702, 27680, 27680, 27680, 27680, 27653, 27653, 27653, 27653, 27653, 27630, 27630, 27630, 27630, 27603, 27603, 27603, 27603, 27581, 27581, 27581, 27581, 27581, 27553, 27553, 27553, 27553, 27531, 27531, 27531, 27531, 27503, 27503, 27503, 27503, 27503, 27481, 27481, 27481, 27481, 27453, 27453, 27453, 27453, 27431, 27431, 27431, 27431, 27431, 27403, 27403, 27403, 27403, 27381, 27381, 27381, 27381, 27353, 27353, 27353, 27353, 27353, 27331, 27331, 27331, 27331, 27303, 27303, 27303, 27303, 27281, 27281, 27281, 27281, 27281, 27253, 27253, 27253, 27253, 27231, 27231, 27231, 27231, 27209, 27209, 27209, 27209, 27209, 27181, 27181, 27181, 27181, 27159, 27159, 27159, 27159, 27159, 27131, 27131, 27131, 27131, 27109, 27109, 27109, 27109, 27081, 27081, 27081, 27081, 27081, 27059, 27059, 27059, 27059, 27031, 27031, 27031, 27031, 27009, 27009, 27009, 27009, 27009, 26981, 26981, 26981, 26981, 26959, 26959, 26959, 26959, 26959, 26931, 26931, 26931, 26931, 26909, 26909, 26909, 26909, 26881, 26881, 26881, 26881, 26881, 26859, 26859, 26859, 26859, 26831, 26831, 26831, 26831, 26831, 26809, 26809, 26809, 26809, 26781, 26781, 26781, 26781, 26759, 26759, 26759, 26759, 26759, 26731, 26731, 26731, 26731, 26709, 26709, 26709, 26709, 26709, 26681, 26681, 26681, 26681, 26659, 26659, 26659, 26659, 26631, 26631, 26631, 26631, 26631, 26609, 26609, 26609, 26609, 26581, 26581, 26581, 26581, 26581, 26559, 26559, 26559, 26559, 26531, 26531, 26531, 26531, 26509, 26509, 26509, 26509, 26509, 26481, 26481, 26481, 26481, 26459, 26459, 26459, 26459, 26459, 26431, 26431, 26431, 26431, 26408, 26408, 26408, 26408, 26408, 26381, 26381, 26381, 26381, 26358, 26358, 26358, 26358, 26330, 26330, 26330, 26330, 26330, 26308, 26308, 26308, 26308, 26280, 26280, 26280, 26280, 26280, 26258, 26258, 26258, 26258, 26230, 26230, 26230, 26230, 26230, 26208, 26208, 26208, 26208, 26180, 26180, 26180, 26180, 26158, 26158, 26158, 26158, 26158, 26130, 26130, 26130, 26130, 26107, 26107, 26107, 26107, 26107, 26085, 26085, 26085, 26085, 26057, 26057, 26057, 26057, 26057, 26035, 26035, 26035, 26035, 26007, 26007, 26007, 26007, 26007, 25985, 25985, 25985, 25985, 25957, 25957, 25957, 25957, 25957, 25934, 25934, 25934, 25934, 25906, 25906, 25906, 25906, 25884, 25884, 25884, 25884, 25884, 25856, 25856, 25856, 25856, 25834, 25834, 25834, 25834, 25834, 25806, 25806, 25806, 25806, 25784, 25784, 25784, 25784, 25784, 25756, 25756, 25756, 25756, 25733, 25733, 25733, 25733, 25733, 25705, 25705, 25705, 25705, 25683, 25683, 25683, 25683, 25683, 25655, 25655, 25655, 25655, 25633, 25633, 25633, 25633, 25633, 25605, 25605, 25605, 25605, 25582, 25582, 25582, 25582, 25582, 25554, 25554, 25554, 25554, 25532, 25532, 25532, 25532, 25532, 25504, 25504, 25504, 25504, 25482, 25482, 25482, 25482, 25482, 25454, 25454, 25454, 25454, 25431, 25431, 25431, 25431, 25431, 25403, 25403, 25403, 25403, 25381, 25381, 25381, 25381, 25381, 25353, 25353, 25353, 25353, 25330, 25330, 25330, 25330, 25330, 25302, 25302, 25302, 25302, 25280, 25280, 25280, 25280, 25280, 25252, 25252, 25252, 25252, 25230, 25230, 25230, 25230, 25230, 25202, 25202, 25202, 25202, 25179, 25179, 25179, 25179, 25179, 25151, 25151, 25151, 25151, 25151, 25129, 25129, 25129, 25129, 25101, 25101, 25101, 25101, 25101, 25078, 25078, 25078, 25078, 25050, 25050, 25050, 25050, 25050, 25028, 25028, 25028, 25028, 25005, 25005, 25005, 25005, 25005, 24977, 24977, 24977, 24977, 24955, 24955, 24955, 24955, 24955, 24927, 24927, 24927, 24927, 24904, 24904, 24904, 24904, 24904, 24876, 24876, 24876, 24876, 24876, 24854, 24854, 24854, 24854, 24826, 24826, 24826, 24826, 24826, 24803, 24803, 24803, 24803, 24775, 24775, 24775, 24775, 24775, 24753, 24753, 24753, 24753, 24725, 24725, 24725, 24725, 24725, 24702, 24702, 24702, 24702, 24702, 24674, 24674, 24674, 24674, 24652, 24652, 24652, 24652, 24652, 24623, 24623, 24623, 24623, 24601, 24601, 24601, 24601, 24601, 24573, 24573, 24573, 24573, 24550, 24550, 24550, 24550, 24550, 24522, 24522, 24522, 24522, 24522, 24500, 24500, 24500, 24500, 24472, 24472, 24472, 24472, 24472, 24449, 24449, 24449, 24449, 24421, 24421, 24421, 24421, 24421, 24398, 24398, 24398, 24398, 24398, 24370, 24370, 24370, 24370, 24348, 24348, 24348, 24348, 24348, 24320, 24320, 24320, 24320, 24297, 24297, 24297, 24297, 24297, 24269, 24269, 24269, 24269, 24269, 24246, 24246, 24246, 24246, 24218, 24218, 24218, 24218, 24218, 24196, 24196, 24196, 24196, 24167, 24167, 24167, 24167, 24167, 24145, 24145, 24145, 24145, 24145, 24117, 24117, 24117, 24117, 24094, 24094, 24094, 24094, 24094, 24066, 24066, 24066, 24066, 24066, 24043, 24043, 24043, 24043, 24015, 24015, 24015, 24015, 24015, 23993, 23993, 23993, 23993, 23993, 23964, 23964, 23964, 23964, 23942, 23942, 23942, 23942, 23942, 23914, 23914, 23914, 23914, 23891, 23891, 23891, 23891, 23891, 23868, 23868, 23868, 23868, 23868, 23840, 23840, 23840, 23840, 23818, 23818, 23818, 23818, 23818, 23789, 23789, 23789, 23789, 23789, 23767, 23767, 23767, 23767, 23738, 23738, 23738, 23738, 23738, 23716, 23716, 23716, 23716, 23716, 23688, 23688, 23688, 23688, 23665, 23665, 23665, 23665, 23665, 23637, 23637, 23637, 23637, 23637, 23614, 23614, 23614, 23614, 23586, 23586, 23586, 23586, 23586, 23563, 23563, 23563, 23563, 23563, 23535, 23535, 23535, 23535, 23512, 23512, 23512, 23512, 23512, 23484, 23484, 23484, 23484, 23484, 23461, 23461, 23461, 23461, 23461, 23433, 23433, 23433, 23433, 23410, 23410, 23410, 23410, 23410, 23382, 23382, 23382, 23382, 23382, 23359, 23359, 23359, 23359, 23331, 23331, 23331, 23331, 23331, 23308, 23308, 23308, 23308, 23308, 23280, 23280, 23280, 23280, 23257, 23257, 23257, 23257, 23257, 23229, 23229, 23229, 23229, 23229, 23206, 23206, 23206, 23206, 23206, 23178, 23178, 23178, 23178, 23155, 23155, 23155, 23155, 23155, 23127, 23127, 23127, 23127, 23127, 23104, 23104, 23104, 23104, 23076, 23076, 23076, 23076, 23076, 23053, 23053, 23053, 23053, 23053, 23025, 23025, 23025, 23025, 23025, 23002, 23002, 23002, 23002, 22974, 22974, 22974, 22974, 22974, 22951, 22951, 22951, 22951, 22951, 22922, 22922, 22922, 22922, 22922, 22900, 22900, 22900, 22900, 22871, 22871, 22871, 22871, 22871, 22849, 22849, 22849, 22849, 22849, 22820, 22820, 22820, 22820, 22820, 22797, 22797, 22797, 22797, 22769, 22769, 22769, 22769, 22769, 22746, 22746, 22746, 22746, 22746, 22724, 22724, 22724, 22724, 22724, 22695, 22695, 22695, 22695, 22672, 22672, 22672, 22672, 22672, 22644, 22644, 22644, 22644, 22644, 22621, 22621, 22621, 22621, 22621, 22593, 22593, 22593, 22593, 22593, 22570, 22570, 22570, 22570, 22541, 22541, 22541, 22541, 22541, 22519, 22519, 22519, 22519, 22519, 22490, 22490, 22490, 22490, 22490, 22467, 22467, 22467, 22467, 22439, 22439, 22439, 22439, 22439, 22416, 22416, 22416, 22416, 22416, 22388, 22388, 22388, 22388, 22388, 22365, 22365, 22365, 22365, 22365, 22336, 22336, 22336, 22336, 22313, 22313, 22313, 22313, 22313, 22285, 22285, 22285, 22285, 22285, 22262, 22262, 22262, 22262, 22262, 22234, 22234, 22234, 22234, 22234, 22211, 22211, 22211, 22211, 22211, 22182, 22182, 22182, 22182, 22159, 22159, 22159, 22159, 22159, 22131, 22131, 22131, 22131, 22131, 22108, 22108, 22108, 22108, 22108, 22079, 22079, 22079, 22079, 22079, 22057, 22057, 22057, 22057, 22057, 22028, 22028, 22028, 22028, 22005, 22005, 22005, 22005, 22005, 21977, 21977, 21977, 21977, 21977, 21954, 21954, 21954, 21954, 21954, 21925, 21925, 21925, 21925, 21925, 21902, 21902, 21902, 21902, 21902, 21874, 21874, 21874, 21874, 21851, 21851, 21851, 21851, 21851, 21822, 21822, 21822, 21822, 21822, 21799, 21799, 21799, 21799, 21799, 21771, 21771, 21771, 21771, 21771, 21748, 21748, 21748, 21748, 21748, 21719, 21719, 21719, 21719, 21719, 21696, 21696, 21696, 21696, 21696, 21668, 21668, 21668, 21668, 21645, 21645, 21645, 21645, 21645, 21616, 21616, 21616, 21616, 21616, 21593, 21593, 21593, 21593, 21593, 21570, 21570, 21570, 21570, 21570, 21541, 21541, 21541, 21541, 21541, 21518, 21518, 21518, 21518, 21518, 21490, 21490, 21490, 21490, 21490, 21467, 21467, 21467, 21467, 21467, 21438, 21438, 21438, 21438, 21415, 21415, 21415, 21415, 21415, 21387, 21387, 21387, 21387, 21387, 21364, 21364, 21364, 21364, 21364, 21335, 21335, 21335, 21335, 21335, 21312, 21312, 21312, 21312, 21312, 21283, 21283, 21283, 21283, 21283, 21260, 21260, 21260, 21260, 21260, 21231, 21231, 21231, 21231, 21231, 21208, 21208, 21208, 21208, 21208, 21180, 21180, 21180, 21180, 21180, 21157, 21157, 21157, 21157, 21157, 21128, 21128, 21128, 21128, 21128, 21105, 21105, 21105, 21105, 21076, 21076, 21076, 21076, 21076, 21053, 21053, 21053, 21053, 21053, 21024, 21024, 21024, 21024, 21024, 21001, 21001, 21001, 21001, 21001, 20973, 20973, 20973, 20973, 20973, 20950, 20950, 20950, 20950, 20950, 20921, 20921, 20921, 20921, 20921, 20898, 20898, 20898, 20898, 20898, 20869, 20869, 20869, 20869, 20869, 20846, 20846, 20846, 20846, 20846, 20817, 20817, 20817, 20817, 20817, 20794, 20794, 20794, 20794, 20794, 20765, 20765, 20765, 20765, 20765, 20742, 20742, 20742, 20742, 20742, 20713, 20713, 20713, 20713, 20713, 20690, 20690, 20690, 20690, 20690, 20661, 20661, 20661, 20661, 20661, 20638, 20638, 20638, 20638, 20638, 20609, 20609, 20609, 20609, 20609, 20586, 20586, 20586, 20586, 20586, 20557, 20557, 20557, 20557, 20557, 20534, 20534, 20534, 20534, 20534, 20505, 20505, 20505, 20505, 20505, 20482, 20482, 20482, 20482, 20482, 20453, 20453, 20453, 20453, 20453, 20430, 20430, 20430, 20430, 20430, 20407, 20407, 20407, 20407, 20407, 20378, 20378, 20378, 20378, 20378, 20355, 20355, 20355, 20355, 20355, 20326, 20326, 20326, 20326, 20326, 20303, 20303, 20303, 20303, 20303, 20274, 20274, 20274, 20274, 20274, 20251, 20251, 20251, 20251, 20251, 20222, 20222, 20222, 20222, 20222, 20199, 20199, 20199, 20199, 20199, 20170, 20170, 20170, 20170, 20170, 20147, 20147, 20147, 20147, 20147, 20147, 20118, 20118, 20118, 20118, 20118, 20095, 20095, 20095, 20095, 20095, 20066, 20066, 20066, 20066, 20066, 20042, 20042, 20042, 20042, 20042, 20013, 20013, 20013, 20013, 20013, 19990, 19990, 19990, 19990, 19990, 19961, 19961, 19961, 19961, 19961, 19938, 19938, 19938, 19938, 19938, 19909, 19909, 19909, 19909, 19909, 19886, 19886, 19886, 19886, 19886, 19857, 19857, 19857, 19857, 19857, 19834, 19834, 19834, 19834, 19834, 19805, 19805, 19805, 19805, 19805, 19805, 19781, 19781, 19781, 19781, 19781, 19752, 19752, 19752, 19752, 19752, 19729, 19729, 19729, 19729, 19729, 19700, 19700, 19700, 19700, 19700, 19677, 19677, 19677, 19677, 19677, 19648, 19648, 19648, 19648, 19648, 19624, 19624, 19624, 19624, 19624, 19595, 19595, 19595, 19595, 19595, 19595, 19572, 19572, 19572, 19572, 19572, 19543, 19543, 19543, 19543, 19543, 19520, 19520, 19520, 19520, 19520, 19490, 19490, 19490, 19490, 19490, 19467, 19467, 19467, 19467, 19467, 19438, 19438, 19438, 19438, 19438, 19415, 19415, 19415, 19415, 19415, 19415, 19386, 19386, 19386, 19386, 19386, 19362, 19362, 19362, 19362, 19362, 19333, 19333, 19333, 19333, 19333, 19310, 19310, 19310, 19310, 19310, 19287, 19287, 19287, 19287, 19287, 19257, 19257, 19257, 19257, 19257, 19257, 19234, 19234, 19234, 19234, 19234, 19205, 19205, 19205, 19205, 19205, 19181, 19181, 19181, 19181, 19181, 19152, 19152, 19152, 19152, 19152, 19129, 19129, 19129, 19129, 19129, 19100, 19100, 19100, 19100, 19100, 19100, 19076, 19076, 19076, 19076, 19076, 19047, 19047, 19047, 19047, 19047, 19024, 19024, 19024, 19024, 19024, 18995, 18995, 18995, 18995, 18995, 18971, 18971, 18971, 18971, 18971, 18971, 18942, 18942, 18942, 18942, 18942, 18919, 18919, 18919, 18919, 18919, 18889, 18889, 18889, 18889, 18889, 18866, 18866, 18866, 18866, 18866, 18866, 18837, 18837, 18837, 18837, 18837, 18813, 18813, 18813, 18813, 18813, 18784, 18784, 18784, 18784, 18784, 18760, 18760, 18760, 18760, 18760, 18760, 18731, 18731, 18731, 18731, 18731, 18708, 18708, 18708, 18708, 18708, 18678, 18678, 18678, 18678, 18678, 18655, 18655, 18655, 18655, 18655, 18655, 18626, 18626, 18626, 18626, 18626, 18602, 18602, 18602, 18602, 18602, 18573, 18573, 18573, 18573, 18573, 18549, 18549, 18549, 18549, 18549, 18549, 18520, 18520, 18520, 18520, 18520, 18497, 18497, 18497, 18497, 18497, 18467, 18467, 18467, 18467, 18467, 18444, 18444, 18444, 18444, 18444, 18444, 18414, 18414, 18414, 18414, 18414, 18391, 18391, 18391, 18391, 18391, 18362, 18362, 18362, 18362, 18362, 18362, 18338, 18338, 18338, 18338, 18338, 18309, 18309, 18309, 18309, 18309, 18285, 18285, 18285, 18285, 18285, 18285, 18256, 18256, 18256, 18256, 18256, 18232, 18232, 18232, 18232, 18232, 18203, 18203, 18203, 18203, 18203, 18179, 18179, 18179, 18179, 18179, 18179, 18150, 18150, 18150, 18150, 18150, 18126, 18126, 18126, 18126, 18126, 18103, 18103, 18103, 18103, 18103, 18103, 18073, 18073, 18073, 18073, 18073, 18050, 18050, 18050, 18050, 18050, 18050, 18020, 18020, 18020, 18020, 18020, 17997, 17997, 17997, 17997, 17997, 17967, 17967, 17967, 17967, 17967, 17967, 17944, 17944, 17944, 17944, 17944, 17914, 17914, 17914, 17914, 17914, 17890, 17890, 17890, 17890, 17890, 17890, 17861, 17861, 17861, 17861, 17861, 17837, 17837, 17837, 17837, 17837, 17808, 17808, 17808, 17808, 17808, 17808, 17784, 17784, 17784, 17784, 17784, 17755, 17755, 17755, 17755, 17755, 17755, 17731, 17731, 17731, 17731, 17731, 17701, 17701, 17701, 17701, 17701, 17678, 17678, 17678, 17678, 17678, 17678, 17648, 17648, 17648, 17648, 17648, 17625, 17625, 17625, 17625, 17625, 17625, 17595, 17595, 17595, 17595, 17595, 17571, 17571, 17571, 17571, 17571, 17542, 17542, 17542, 17542, 17542, 17542, 17518, 17518, 17518, 17518, 17518, 17489, 17489, 17489, 17489, 17489, 17489, 17465, 17465, 17465, 17465, 17465, 17435, 17435, 17435, 17435, 17435, 17435, 17412, 17412, 17412, 17412, 17412, 17382, 17382, 17382, 17382, 17382, 17358, 17358, 17358, 17358, 17358, 17358, 17329, 17329, 17329, 17329, 17329, 17305, 17305, 17305, 17305, 17305, 17305, 17275, 17275, 17275, 17275, 17275, 17251, 17251, 17251, 17251, 17251, 17251, 17222, 17222, 17222, 17222, 17222, 17198, 17198, 17198, 17198, 17198, 17198, 17168, 17168, 17168, 17168, 17168, 17145, 17145, 17145, 17145, 17145, 17145, 17115, 17115, 17115, 17115, 17115, 17091, 17091, 17091, 17091, 17091, 17091, 17061, 17061, 17061, 17061, 17061, 17038, 17038, 17038, 17038, 17038, 17038, 17008, 17008, 17008, 17008, 17008, 16984, 16984, 16984, 16984, 16984, 16984, 16954, 16954, 16954, 16954, 16954, 16931, 16931, 16931, 16931, 16931, 16931, 16907, 16907, 16907, 16907, 16907, 16877, 16877, 16877, 16877, 16877, 16877, 16853, 16853, 16853, 16853, 16853, 16823, 16823, 16823, 16823, 16823, 16823, 16800, 16800, 16800, 16800, 16800, 16770, 16770, 16770, 16770, 16770, 16770, 16746, 16746, 16746, 16746, 16746, 16716, 16716, 16716, 16716, 16716, 16716, 16692, 16692, 16692, 16692, 16692, 16692, 16662, 16662, 16662, 16662, 16662, 16639, 16639, 16639, 16639, 16639, 16639, 16609, 16609, 16609, 16609, 16609, 16585, 16585, 16585, 16585, 16585, 16585, 16555, 16555, 16555, 16555, 16555, 16531, 16531, 16531, 16531, 16531, 16531, 16501, 16501, 16501, 16501, 16501, 16501, 16477, 16477, 16477, 16477, 16477, 16448, 16448, 16448, 16448, 16448, 16448, 16424, 16424, 16424, 16424, 16424, 16394, 16394, 16394, 16394, 16394, 16394, 16370, 16370, 16370, 16370, 16370, 16370, 16340, 16340, 16340, 16340, 16340, 16316, 16316, 16316, 16316, 16316, 16316, 16286, 16286, 16286, 16286, 16286, 16286, 16262, 16262, 16262, 16262, 16262, 16232, 16232, 16232, 16232, 16232, 16232, 16208, 16208, 16208, 16208, 16208, 16178, 16178, 16178, 16178, 16178, 16178, 16154, 16154, 16154, 16154, 16154, 16154, 16124, 16124, 16124, 16124, 16124, 16100, 16100, 16100, 16100, 16100, 16100, 16070, 16070, 16070, 16070, 16070, 16070, 16046, 16046, 16046, 16046, 16046, 16016, 16016, 16016, 16016, 16016, 16016, 15992, 15992, 15992, 15992, 15992, 15992, 15962, 15962, 15962, 15962, 15962, 15938, 15938, 15938, 15938, 15938, 15938, 15908, 15908, 15908, 15908, 15908, 15908, 15884, 15884, 15884, 15884, 15884, 15884, 15854, 15854, 15854, 15854, 15854, 15830, 15830, 15830, 15830, 15830, 15830, 15800, 15800, 15800, 15800, 15800, 15800, 15776, 15776, 15776, 15776, 15776, 15746, 15746, 15746, 15746, 15746, 15746, 15722, 15722, 15722, 15722, 15722, 15722, 15698, 15698, 15698, 15698, 15698, 15698, 15668, 15668, 15668, 15668, 15668, 15644, 15644, 15644, 15644, 15644, 15644, 15614, 15614, 15614, 15614, 15614, 15614, 15590, 15590, 15590, 15590, 15590, 15590, 15559, 15559, 15559, 15559, 15559, 15535, 15535, 15535, 15535, 15535, 15535, 15505, 15505, 15505, 15505, 15505, 15505, 15481, 15481, 15481, 15481, 15481, 15481, 15451, 15451, 15451, 15451, 15451, 15427, 15427, 15427, 15427, 15427, 15427, 15397, 15397, 15397, 15397, 15397, 15397, 15372, 15372, 15372, 15372, 15372, 15372, 15342, 15342, 15342, 15342, 15342, 15342, 15318, 15318, 15318, 15318, 15318, 15288, 15288, 15288, 15288, 15288, 15288, 15264, 15264, 15264, 15264, 15264, 15264, 15233, 15233, 15233, 15233, 15233, 15233, 15209, 15209, 15209, 15209, 15209, 15209, 15179, 15179, 15179, 15179, 15179, 15179, 15155, 15155, 15155, 15155, 15155, 15125, 15125, 15125, 15125, 15125, 15125, 15100, 15100, 15100, 15100, 15100, 15100, 15070, 15070, 15070, 15070, 15070, 15070, 15046, 15046, 15046, 15046, 15046, 15046, 15016, 15016, 15016, 15016, 15016, 15016, 14991, 14991, 14991, 14991, 14991, 14991, 14961, 14961, 14961, 14961, 14961, 14937, 14937, 14937, 14937, 14937, 14937, 14907, 14907, 14907, 14907, 14907, 14907, 14882, 14882, 14882, 14882, 14882, 14882, 14852, 14852, 14852, 14852, 14852, 14852, 14828, 14828, 14828, 14828, 14828, 14828, 14797, 14797, 14797, 14797, 14797, 14797, 14773, 14773, 14773, 14773, 14773, 14773, 14743, 14743, 14743, 14743, 14743, 14743, 14718, 14718, 14718, 14718, 14718, 14718, 14688, 14688, 14688, 14688, 14688, 14688, 14664, 14664, 14664, 14664, 14664, 14633, 14633, 14633, 14633, 14633, 14633, 14609, 14609, 14609, 14609, 14609, 14609, 14579, 14579, 14579, 14579, 14579, 14579, 14554, 14554, 14554, 14554, 14554, 14554, 14530, 14530, 14530, 14530, 14530, 14530, 14499, 14499, 14499, 14499, 14499, 14499, 14475, 14475, 14475, 14475, 14475, 14475, 14445, 14445, 14445, 14445, 14445, 14445, 14420, 14420, 14420, 14420, 14420, 14420, 14390, 14390, 14390, 14390, 14390, 14390, 14365, 14365, 14365, 14365, 14365, 14365, 14335, 14335, 14335, 14335, 14335, 14335, 14311, 14311, 14311, 14311, 14311, 14311, 14280, 14280, 14280, 14280, 14280, 14280, 14256, 14256, 14256, 14256, 14256, 14256, 14225, 14225, 14225, 14225, 14225, 14225, 14201, 14201, 14201, 14201, 14201, 14201, 14170, 14170, 14170, 14170, 14170, 14170, 14146, 14146, 14146, 14146, 14146, 14146, 14115, 14115, 14115, 14115, 14115, 14115, 14091, 14091, 14091, 14091, 14091, 14091, 14060, 14060, 14060, 14060, 14060, 14060, 14060, 14036, 14036, 14036, 14036, 14036, 14036, 14005, 14005, 14005, 14005, 14005, 14005, 13981, 13981, 13981, 13981, 13981, 13981, 13950, 13950, 13950, 13950, 13950, 13950, 13925, 13925, 13925, 13925, 13925, 13925, 13895, 13895, 13895, 13895, 13895, 13895, 13870, 13870, 13870, 13870, 13870, 13870, 13840, 13840, 13840, 13840, 13840, 13840, 13815, 13815, 13815, 13815, 13815, 13815, 13785, 13785, 13785, 13785, 13785, 13785, 13785, 13760, 13760, 13760, 13760, 13760, 13760, 13729, 13729, 13729, 13729, 13729, 13729, 13705, 13705, 13705, 13705, 13705, 13705, 13674, 13674, 13674, 13674, 13674, 13674, 13650, 13650, 13650, 13650, 13650, 13650, 13619, 13619, 13619, 13619, 13619, 13619, 13594, 13594, 13594, 13594, 13594, 13594, 13594, 13564, 13564, 13564, 13564, 13564, 13564, 13539, 13539, 13539, 13539, 13539, 13539, 13508, 13508, 13508, 13508, 13508, 13508, 13484, 13484, 13484, 13484, 13484, 13484, 13453, 13453, 13453, 13453, 13453, 13453, 13453, 13428, 13428, 13428, 13428, 13428, 13428, 13397, 13397, 13397, 13397, 13397, 13397, 13373, 13373, 13373, 13373, 13373, 13373, 13342, 13342, 13342, 13342, 13342, 13342, 13317, 13317, 13317, 13317, 13317, 13317, 13317, 13293, 13293, 13293, 13293, 13293, 13293, 13262, 13262, 13262, 13262, 13262, 13262, 13237, 13237, 13237, 13237, 13237, 13237, 13206, 13206, 13206, 13206, 13206, 13206, 13206, 13182, 13182, 13182, 13182, 13182, 13182, 13151, 13151, 13151, 13151, 13151, 13151, 13126, 13126, 13126, 13126, 13126, 13126, 13095, 13095, 13095, 13095, 13095, 13095, 13095, 13071, 13071, 13071, 13071, 13071, 13071, 13040, 13040, 13040, 13040, 13040, 13040, 13015, 13015, 13015, 13015, 13015, 13015, 13015, 12984, 12984, 12984, 12984, 12984, 12984, 12959, 12959, 12959, 12959, 12959, 12959, 12928, 12928, 12928, 12928, 12928, 12928, 12928, 12904, 12904, 12904, 12904, 12904, 12904, 12873, 12873, 12873, 12873, 12873, 12873, 12848, 12848, 12848, 12848, 12848, 12848, 12848, 12817, 12817, 12817, 12817, 12817, 12817, 12792, 12792, 12792, 12792, 12792, 12792, 12761, 12761, 12761, 12761, 12761, 12761, 12761, 12736, 12736, 12736, 12736, 12736, 12736, 12705, 12705, 12705, 12705, 12705, 12705, 12705, 12681, 12681, 12681, 12681, 12681, 12681, 12650, 12650, 12650, 12650, 12650, 12650, 12625, 12625, 12625, 12625, 12625, 12625, 12625, 12594, 12594, 12594, 12594, 12594, 12594, 12569, 12569, 12569, 12569, 12569, 12569, 12569, 12538, 12538, 12538, 12538, 12538, 12538, 12513, 12513, 12513, 12513, 12513, 12513, 12482, 12482, 12482, 12482, 12482, 12482, 12482, 12457, 12457, 12457, 12457, 12457, 12457, 12426, 12426, 12426, 12426, 12426, 12426, 12426, 12401, 12401, 12401, 12401, 12401, 12401, 12370, 12370, 12370, 12370, 12370, 12370, 12370, 12345, 12345, 12345, 12345, 12345, 12345, 12314, 12314, 12314, 12314, 12314, 12314, 12314, 12289, 12289, 12289, 12289, 12289, 12289, 12258, 12258, 12258, 12258, 12258, 12258, 12258, 12233, 12233, 12233, 12233, 12233, 12233, 12202, 12202, 12202, 12202, 12202, 12202, 12202, 12177, 12177, 12177, 12177, 12177, 12177, 12146, 12146, 12146, 12146, 12146, 12146, 12146, 12121, 12121, 12121, 12121, 12121, 12121, 12090, 12090, 12090, 12090, 12090, 12090, 12090, 12065, 12065, 12065, 12065, 12065, 12065, 12040, 12040, 12040, 12040, 12040, 12040, 12040, 12008, 12008, 12008, 12008, 12008, 12008, 12008, 11983, 11983, 11983, 11983, 11983, 11983, 11952, 11952, 11952, 11952, 11952, 11952, 11952, 11927, 11927, 11927, 11927, 11927, 11927, 11896, 11896, 11896, 11896, 11896, 11896, 11896, 11871, 11871, 11871, 11871, 11871, 11871, 11871, 11840, 11840, 11840, 11840, 11840, 11840, 11815, 11815, 11815, 11815, 11815, 11815, 11815, 11783, 11783, 11783, 11783, 11783, 11783, 11758, 11758, 11758, 11758, 11758, 11758, 11758, 11727, 11727, 11727, 11727, 11727, 11727, 11727, 11702, 11702, 11702, 11702, 11702, 11702, 11670, 11670, 11670, 11670, 11670, 11670, 11670, 11645, 11645, 11645, 11645, 11645, 11645, 11645, 11614, 11614, 11614, 11614, 11614, 11614, 11589, 11589, 11589, 11589, 11589, 11589, 11589, 11558, 11558, 11558, 11558, 11558, 11558, 11558, 11532, 11532, 11532, 11532, 11532, 11532, 11501, 11501, 11501, 11501, 11501, 11501, 11501, 11476, 11476, 11476, 11476, 11476, 11476, 11476, 11444, 11444, 11444, 11444, 11444, 11444, 11444, 11419, 11419, 11419, 11419, 11419, 11419, 11388, 11388, 11388, 11388, 11388, 11388, 11388, 11363, 11363, 11363, 11363, 11363, 11363, 11363, 11331, 11331, 11331, 11331, 11331, 11331, 11331, 11306, 11306, 11306, 11306, 11306, 11306, 11275, 11275, 11275, 11275, 11275, 11275, 11275, 11249, 11249, 11249, 11249, 11249, 11249, 11249, 11218, 11218, 11218, 11218, 11218, 11218, 11218, 11193, 11193, 11193, 11193, 11193, 11193, 11193, 11161, 11161, 11161, 11161, 11161, 11161, 11136, 11136, 11136, 11136, 11136, 11136, 11136, 11104, 11104, 11104, 11104, 11104, 11104, 11104, 11079, 11079, 11079, 11079, 11079, 11079, 11079, 11048, 11048, 11048, 11048, 11048, 11048, 11048, 11022, 11022, 11022, 11022, 11022, 11022, 11022, 10991, 10991, 10991, 10991, 10991, 10991, 10991, 10966, 10966, 10966, 10966, 10966, 10966, 10934, 10934, 10934, 10934, 10934, 10934, 10934, 10909, 10909, 10909, 10909, 10909, 10909, 10909, 10877, 10877, 10877, 10877, 10877, 10877, 10877, 10852, 10852, 10852, 10852, 10852, 10852, 10852, 10820, 10820, 10820, 10820, 10820, 10820, 10820, 10795, 10795, 10795, 10795, 10795, 10795, 10795, 10769, 10769, 10769, 10769, 10769, 10769, 10769, 10738, 10738, 10738, 10738, 10738, 10738, 10738, 10712, 10712, 10712, 10712, 10712, 10712, 10712, 10681, 10681, 10681, 10681, 10681, 10681, 10681, 10655, 10655, 10655, 10655, 10655, 10655, 10655, 10624, 10624, 10624, 10624, 10624, 10624, 10624, 10598, 10598, 10598, 10598, 10598, 10598, 10598, 10567, 10567, 10567, 10567, 10567, 10567, 10567, 10541, 10541, 10541, 10541, 10541, 10541, 10541, 10509, 10509, 10509, 10509, 10509, 10509, 10509, 10484, 10484, 10484, 10484, 10484, 10484, 10484, 10452, 10452, 10452, 10452, 10452, 10452, 10452, 10427, 10427, 10427, 10427, 10427, 10427, 10427, 10395, 10395, 10395, 10395, 10395, 10395, 10395, 10370, 10370, 10370, 10370, 10370, 10370, 10370, 10338, 10338, 10338, 10338, 10338, 10338, 10338, 10312, 10312, 10312, 10312, 10312, 10312, 10312, 10281, 10281, 10281, 10281, 10281, 10281, 10281, 10255, 10255, 10255, 10255, 10255, 10255, 10255, 10255, 10223, 10223, 10223, 10223, 10223, 10223, 10223, 10198, 10198, 10198, 10198, 10198, 10198, 10198, 10166, 10166, 10166, 10166, 10166, 10166, 10166, 10140, 10140, 10140, 10140, 10140, 10140, 10140, 10108, 10108, 10108, 10108, 10108, 10108, 10108, 10083, 10083, 10083, 10083, 10083, 10083, 10083, 10051, 10051, 10051, 10051, 10051, 10051, 10051, 10051, 10025, 10025, 10025, 10025, 10025, 10025, 10025, 9994, 9994, 9994, 9994, 9994, 9994, 9994, 9968, 9968, 9968, 9968, 9968, 9968, 9968, 9936, 9936, 9936, 9936, 9936, 9936, 9936, 9936, 9910, 9910, 9910, 9910, 9910, 9910, 9910, 9878, 9878, 9878, 9878, 9878, 9878, 9878, 9853, 9853, 9853, 9853, 9853, 9853, 9853, 9821, 9821, 9821, 9821, 9821, 9821, 9821, 9821, 9795, 9795, 9795, 9795, 9795, 9795, 9795, 9763, 9763, 9763, 9763, 9763, 9763, 9763, 9738, 9738, 9738, 9738, 9738, 9738, 9738, 9738, 9706, 9706, 9706, 9706, 9706, 9706, 9706, 9680, 9680, 9680, 9680, 9680, 9680, 9680, 9648, 9648, 9648, 9648, 9648, 9648, 9648, 9648, 9622, 9622, 9622, 9622, 9622, 9622, 9622, 9590, 9590, 9590, 9590, 9590, 9590, 9590, 9564, 9564, 9564, 9564, 9564, 9564, 9564, 9564, 9532, 9532, 9532, 9532, 9532, 9532, 9532, 9507, 9507, 9507, 9507, 9507, 9507, 9507, 9481, 9481, 9481, 9481, 9481, 9481, 9481, 9481, 9449, 9449, 9449, 9449, 9449, 9449, 9449, 9423, 9423, 9423, 9423, 9423, 9423, 9423, 9423, 9391, 9391, 9391, 9391, 9391, 9391, 9391, 9365, 9365, 9365, 9365, 9365, 9365, 9365, 9365, 9333, 9333, 9333, 9333, 9333, 9333, 9333, 9307, 9307, 9307, 9307, 9307, 9307, 9307, 9307, 9275, 9275, 9275, 9275, 9275, 9275, 9275, 9249, 9249, 9249, 9249, 9249, 9249, 9249, 9249, 9217, 9217, 9217, 9217, 9217, 9217, 9217, 9191, 9191, 9191, 9191, 9191, 9191, 9191, 9191, 9159, 9159, 9159, 9159, 9159, 9159, 9159, 9133, 9133, 9133, 9133, 9133, 9133, 9133, 9133, 9101, 9101, 9101, 9101, 9101, 9101, 9101, 9075, 9075, 9075, 9075, 9075, 9075, 9075, 9075, 9043, 9043, 9043, 9043, 9043, 9043, 9043, 9017, 9017, 9017, 9017, 9017, 9017, 9017, 9017, 8985, 8985, 8985, 8985, 8985, 8985, 8985, 8985, 8959, 8959, 8959, 8959, 8959, 8959, 8959, 8927, 8927, 8927, 8927, 8927, 8927, 8927, 8927, 8901, 8901, 8901, 8901, 8901, 8901, 8901, 8901, 8868, 8868, 8868, 8868, 8868, 8868, 8868, 8842, 8842, 8842, 8842, 8842, 8842, 8842, 8842, 8810, 8810, 8810, 8810, 8810, 8810, 8810, 8810, 8784, 8784, 8784, 8784, 8784, 8784, 8784, 8752, 8752, 8752, 8752, 8752, 8752, 8752, 8752, 8726, 8726, 8726, 8726, 8726, 8726, 8726, 8726, 8693, 8693, 8693, 8693, 8693, 8693, 8693, 8668, 8668, 8668, 8668, 8668, 8668, 8668, 8668, 8635, 8635, 8635, 8635, 8635, 8635, 8635, 8635, 8609, 8609, 8609, 8609, 8609, 8609, 8609, 8609, 8577, 8577, 8577, 8577, 8577, 8577, 8577, 8577, 8551, 8551, 8551, 8551, 8551, 8551, 8551, 8518, 8518, 8518, 8518, 8518, 8518, 8518, 8518, 8492, 8492, 8492, 8492, 8492, 8492, 8492, 8492, 8460, 8460, 8460, 8460, 8460, 8460, 8460, 8460, 8434, 8434, 8434, 8434, 8434, 8434, 8434, 8434, 8401, 8401, 8401, 8401, 8401, 8401, 8401, 8401, 8375, 8375, 8375, 8375, 8375, 8375, 8375, 8375, 8343, 8343, 8343, 8343, 8343, 8343, 8343, 8316, 8316, 8316, 8316, 8316, 8316, 8316, 8316, 8284, 8284, 8284, 8284, 8284, 8284, 8284, 8284, 8258, 8258, 8258, 8258, 8258, 8258, 8258, 8258, 8232, 8232, 8232, 8232, 8232, 8232, 8232, 8232, 8199, 8199, 8199, 8199, 8199, 8199, 8199, 8199, 8173, 8173, 8173, 8173, 8173, 8173, 8173, 8173, 8140, 8140, 8140, 8140, 8140, 8140, 8140, 8140, 8114, 8114, 8114, 8114, 8114, 8114, 8114, 8114, 8082, 8082, 8082, 8082, 8082, 8082, 8082, 8082, 8056, 8056, 8056, 8056, 8056, 8056, 8056, 8056, 8023, 8023, 8023, 8023, 8023, 8023, 8023, 8023, 7997, 7997, 7997, 7997, 7997, 7997, 7997, 7997, 7964, 7964, 7964, 7964, 7964, 7964, 7964, 7964, 7964, 7938, 7938, 7938, 7938, 7938, 7938, 7938, 7938, 7905, 7905, 7905, 7905, 7905, 7905, 7905, 7905, 7879, 7879, 7879, 7879, 7879, 7879, 7879, 7879, 7846, 7846, 7846, 7846, 7846, 7846, 7846, 7846, 7820, 7820, 7820, 7820, 7820, 7820, 7820, 7820, 7787, 7787, 7787, 7787, 7787, 7787, 7787, 7787, 7761, 7761, 7761, 7761, 7761, 7761, 7761, 7761, 7761, 7728, 7728, 7728, 7728, 7728, 7728, 7728, 7728, 7702, 7702, 7702, 7702, 7702, 7702, 7702, 7702, 7669, 7669, 7669, 7669, 7669, 7669, 7669, 7669, 7643, 7643, 7643, 7643, 7643, 7643, 7643, 7643, 7643, 7610, 7610, 7610, 7610, 7610, 7610, 7610, 7610, 7584, 7584, 7584, 7584, 7584, 7584, 7584, 7584, 7551, 7551, 7551, 7551, 7551, 7551, 7551, 7551, 7551, 7525, 7525, 7525, 7525, 7525, 7525, 7525, 7525, 7492, 7492, 7492, 7492, 7492, 7492, 7492, 7492, 7465, 7465, 7465, 7465, 7465, 7465, 7465, 7465, 7465, 7432, 7432, 7432, 7432, 7432, 7432, 7432, 7432, 7406, 7406, 7406, 7406, 7406, 7406, 7406, 7406, 7373, 7373, 7373, 7373, 7373, 7373, 7373, 7373, 7373, 7347, 7347, 7347, 7347, 7347, 7347, 7347, 7347, 7314, 7314, 7314, 7314, 7314, 7314, 7314, 7314, 7314, 7287, 7287, 7287, 7287, 7287, 7287, 7287, 7287, 7254, 7254, 7254, 7254, 7254, 7254, 7254, 7254, 7254, 7228, 7228, 7228, 7228, 7228, 7228, 7228, 7228, 7195, 7195, 7195, 7195, 7195, 7195, 7195, 7195, 7195, 7169, 7169, 7169, 7169, 7169, 7169, 7169, 7169, 7136, 7136, 7136, 7136, 7136, 7136, 7136, 7136, 7136, 7109, 7109, 7109, 7109, 7109, 7109, 7109, 7109, 7076, 7076, 7076, 7076, 7076, 7076, 7076, 7076, 7076, 7050, 7050, 7050, 7050, 7050, 7050, 7050, 7050, 7050, 7017, 7017, 7017, 7017, 7017, 7017, 7017, 7017, 6990, 6990, 6990, 6990, 6990, 6990, 6990, 6990, 6990, 6957, 6957, 6957, 6957, 6957, 6957, 6957, 6957, 6957, 6931, 6931, 6931, 6931, 6931, 6931, 6931, 6931, 6904, 6904, 6904, 6904, 6904, 6904, 6904, 6904, 6904, 6871, 6871, 6871, 6871, 6871, 6871, 6871, 6871, 6871, 6844, 6844, 6844, 6844, 6844, 6844, 6844, 6844, 6811, 6811, 6811, 6811, 6811, 6811, 6811, 6811, 6811, 6785, 6785, 6785, 6785, 6785, 6785, 6785, 6785, 6785, 6752, 6752, 6752, 6752, 6752, 6752, 6752, 6752, 6752, 6725, 6725, 6725, 6725, 6725, 6725, 6725, 6725, 6725, 6692, 6692, 6692, 6692, 6692, 6692, 6692, 6692, 6692, 6665, 6665, 6665, 6665, 6665, 6665, 6665, 6665, 6632, 6632, 6632, 6632, 6632, 6632, 6632, 6632, 6632, 6605, 6605, 6605, 6605, 6605, 6605, 6605, 6605, 6605, 6572, 6572, 6572, 6572, 6572, 6572, 6572, 6572, 6572, 6545, 6545, 6545, 6545, 6545, 6545, 6545, 6545, 6545, 6512, 6512, 6512, 6512, 6512, 6512, 6512, 6512, 6512, 6486, 6486, 6486, 6486, 6486, 6486, 6486, 6486, 6486, 6452, 6452, 6452, 6452, 6452, 6452, 6452, 6452, 6452, 6426, 6426, 6426, 6426, 6426, 6426, 6426, 6426, 6426, 6392, 6392, 6392, 6392, 6392, 6392, 6392, 6392, 6392, 6366, 6366, 6366, 6366, 6366, 6366, 6366, 6366, 6366, 6332, 6332, 6332, 6332, 6332, 6332, 6332, 6332, 6332, 6305, 6305, 6305, 6305, 6305, 6305, 6305, 6305, 6305, 6272, 6272, 6272, 6272, 6272, 6272, 6272, 6272, 6272, 6272, 6245, 6245, 6245, 6245, 6245, 6245, 6245, 6245, 6245, 6212, 6212, 6212, 6212, 6212, 6212, 6212, 6212, 6212, 6185, 6185, 6185, 6185, 6185, 6185, 6185, 6185, 6185, 6152, 6152, 6152, 6152, 6152, 6152, 6152, 6152, 6152, 6125, 6125, 6125, 6125, 6125, 6125, 6125, 6125, 6125, 6125, 6092, 6092, 6092, 6092, 6092, 6092, 6092, 6092, 6092, 6065, 6065, 6065, 6065, 6065, 6065, 6065, 6065, 6065, 6031, 6031, 6031, 6031, 6031, 6031, 6031, 6031, 6031, 6005, 6005, 6005, 6005, 6005, 6005, 6005, 6005, 6005, 6005, 5971, 5971, 5971, 5971, 5971, 5971, 5971, 5971, 5971, 5944, 5944, 5944, 5944, 5944, 5944, 5944, 5944, 5944, 5944, 5911, 5911, 5911, 5911, 5911, 5911, 5911, 5911, 5911, 5884, 5884, 5884, 5884, 5884, 5884, 5884, 5884, 5884, 5850, 5850, 5850, 5850, 5850, 5850, 5850, 5850, 5850, 5850, 5823, 5823, 5823, 5823, 5823, 5823, 5823, 5823, 5823, 5790, 5790, 5790, 5790, 5790, 5790, 5790, 5790, 5790, 5790, 5763, 5763, 5763, 5763, 5763, 5763, 5763, 5763, 5763, 5729, 5729, 5729, 5729, 5729, 5729, 5729, 5729, 5729, 5729, 5702, 5702, 5702, 5702, 5702, 5702, 5702, 5702, 5702, 5702, 5669, 5669, 5669, 5669, 5669, 5669, 5669, 5669, 5669, 5642, 5642, 5642, 5642, 5642, 5642, 5642, 5642, 5642, 5642, 5608, 5608, 5608, 5608, 5608, 5608, 5608, 5608, 5608, 5608, 5581, 5581, 5581, 5581, 5581, 5581, 5581, 5581, 5581, 5554, 5554, 5554, 5554, 5554, 5554, 5554, 5554, 5554, 5554, 5521, 5521, 5521, 5521, 5521, 5521, 5521, 5521, 5521, 5521, 5494, 5494, 5494, 5494, 5494, 5494, 5494, 5494, 5494, 5494, 5460, 5460, 5460, 5460, 5460, 5460, 5460, 5460, 5460, 5433, 5433, 5433, 5433, 5433, 5433, 5433, 5433, 5433, 5433, 5399, 5399, 5399, 5399, 5399, 5399, 5399, 5399, 5399, 5399, 5372, 5372, 5372, 5372, 5372, 5372, 5372, 5372, 5372, 5372, 5338, 5338, 5338, 5338, 5338, 5338, 5338, 5338, 5338, 5338, 5311, 5311, 5311, 5311, 5311, 5311, 5311, 5311, 5311, 5311, 5278, 5278, 5278, 5278, 5278, 5278, 5278, 5278, 5278, 5278, 5250, 5250, 5250, 5250, 5250, 5250, 5250, 5250, 5250, 5250, 5217, 5217, 5217, 5217, 5217, 5217, 5217, 5217, 5217, 5217, 5190, 5190, 5190, 5190, 5190, 5190, 5190, 5190, 5190, 5190, 5156, 5156, 5156, 5156, 5156, 5156, 5156, 5156, 5156, 5156, 5129, 5129, 5129, 5129, 5129, 5129, 5129, 5129, 5129, 5129, 5095, 5095, 5095, 5095, 5095, 5095, 5095, 5095, 5095, 5095, 5068, 5068, 5068, 5068, 5068, 5068, 5068, 5068, 5068, 5068, 5034, 5034, 5034, 5034, 5034, 5034, 5034, 5034, 5034, 5034, 5034, 5007, 5007, 5007, 5007, 5007, 5007, 5007, 5007, 5007, 5007, 4973, 4973, 4973, 4973, 4973, 4973, 4973, 4973, 4973, 4973, 4945, 4945, 4945, 4945, 4945, 4945, 4945, 4945, 4945, 4945, 4945, 4912, 4912, 4912, 4912, 4912, 4912, 4912, 4912, 4912, 4912, 4884, 4884, 4884, 4884, 4884, 4884, 4884, 4884, 4884, 4884, 4850, 4850, 4850, 4850, 4850, 4850, 4850, 4850, 4850, 4850, 4850, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4789, 4789, 4789, 4789, 4789, 4789, 4789, 4789, 4789, 4789, 4789, 4762, 4762, 4762, 4762, 4762, 4762, 4762, 4762, 4762, 4762, 4728, 4728, 4728, 4728, 4728, 4728, 4728, 4728, 4728, 4728, 4728, 4701, 4701, 4701, 4701, 4701, 4701, 4701, 4701, 4701, 4701, 4667, 4667, 4667, 4667, 4667, 4667, 4667, 4667, 4667, 4667, 4667, 4639, 4639, 4639, 4639, 4639, 4639, 4639, 4639, 4639, 4639, 4605, 4605, 4605, 4605, 4605, 4605, 4605, 4605, 4605, 4605, 4605, 4578, 4578, 4578, 4578, 4578, 4578, 4578, 4578, 4578, 4578, 4578, 4544, 4544, 4544, 4544, 4544, 4544, 4544, 4544, 4544, 4544, 4544, 4516, 4516, 4516, 4516, 4516, 4516, 4516, 4516, 4516, 4516, 4482, 4482, 4482, 4482, 4482, 4482, 4482, 4482, 4482, 4482, 4482, 4455, 4455, 4455, 4455, 4455, 4455, 4455, 4455, 4455, 4455, 4455, 4421, 4421, 4421, 4421, 4421, 4421, 4421, 4421, 4421, 4421, 4421, 4393, 4393, 4393, 4393, 4393, 4393, 4393, 4393, 4393, 4393, 4393, 4359, 4359, 4359, 4359, 4359, 4359, 4359, 4359, 4359, 4359, 4359, 4332, 4332, 4332, 4332, 4332, 4332, 4332, 4332, 4332, 4332, 4332, 4298, 4298, 4298, 4298, 4298, 4298, 4298, 4298, 4298, 4298, 4298, 4270, 4270, 4270, 4270, 4270, 4270, 4270, 4270, 4270, 4270, 4270, 4236, 4236, 4236, 4236, 4236, 4236, 4236, 4236, 4236, 4236, 4236, 4209, 4209, 4209, 4209, 4209, 4209, 4209, 4209, 4209, 4209, 4209, 4209, 4181, 4181, 4181, 4181, 4181, 4181, 4181, 4181, 4181, 4181, 4181, 4147, 4147, 4147, 4147, 4147, 4147, 4147, 4147, 4147, 4147, 4147, 4119, 4119, 4119, 4119, 4119, 4119, 4119, 4119, 4119, 4119, 4119, 4085, 4085, 4085, 4085, 4085, 4085, 4085, 4085, 4085, 4085, 4085, 4085, 4058, 4058, 4058, 4058, 4058, 4058, 4058, 4058, 4058, 4058, 4058, 4023, 4023, 4023, 4023, 4023, 4023, 4023, 4023, 4023, 4023, 4023, 4023, 3996, 3996, 3996, 3996, 3996, 3996, 3996, 3996, 3996, 3996, 3996, 3961, 3961, 3961, 3961, 3961, 3961, 3961, 3961, 3961, 3961, 3961, 3961, 3934, 3934, 3934, 3934, 3934, 3934, 3934, 3934, 3934, 3934, 3934, 3899, 3899, 3899, 3899, 3899, 3899, 3899, 3899, 3899, 3899, 3899, 3899, 3872, 3872, 3872, 3872, 3872, 3872, 3872, 3872, 3872, 3872, 3872, 3837, 3837, 3837, 3837, 3837, 3837, 3837, 3837, 3837, 3837, 3837, 3837, 3810, 3810, 3810, 3810, 3810, 3810, 3810, 3810, 3810, 3810, 3810, 3810, 3775, 3775, 3775, 3775, 3775, 3775, 3775, 3775, 3775, 3775, 3775, 3775, 3748, 3748, 3748, 3748, 3748, 3748, 3748, 3748, 3748, 3748, 3748, 3748, 3713, 3713, 3713, 3713, 3713, 3713, 3713, 3713, 3713, 3713, 3713, 3713, 3686, 3686, 3686, 3686, 3686, 3686, 3686, 3686, 3686, 3686, 3686, 3686, 3651, 3651, 3651, 3651, 3651, 3651, 3651, 3651, 3651, 3651, 3651, 3651, 3624, 3624, 3624, 3624, 3624, 3624, 3624, 3624, 3624, 3624, 3624, 3624, 3589, 3589, 3589, 3589, 3589, 3589, 3589, 3589, 3589, 3589, 3589, 3589, 3561, 3561, 3561, 3561, 3561, 3561, 3561, 3561, 3561, 3561, 3561, 3561, 3527, 3527, 3527, 3527, 3527, 3527, 3527, 3527, 3527, 3527, 3527, 3527, 3499, 3499, 3499, 3499, 3499, 3499, 3499, 3499, 3499, 3499, 3499, 3499, 3465, 3465, 3465, 3465, 3465, 3465, 3465, 3465, 3465, 3465, 3465, 3465, 3465, 3437, 3437, 3437, 3437, 3437, 3437, 3437, 3437, 3437, 3437, 3437, 3437, 3402, 3402, 3402, 3402, 3402, 3402, 3402, 3402, 3402, 3402, 3402, 3402, 3402, 3374, 3374, 3374, 3374, 3374, 3374, 3374, 3374, 3374, 3374, 3374, 3374, 3340, 3340, 3340, 3340, 3340, 3340, 3340, 3340, 3340, 3340, 3340, 3340, 3340, 3312, 3312, 3312, 3312, 3312, 3312, 3312, 3312, 3312, 3312, 3312, 3312, 3277, 3277, 3277, 3277, 3277, 3277, 3277, 3277, 3277, 3277, 3277, 3277, 3277, 3250, 3250, 3250, 3250, 3250, 3250, 3250, 3250, 3250, 3250, 3250, 3250, 3250, 3215, 3215, 3215, 3215, 3215, 3215, 3215, 3215, 3215, 3215, 3215, 3215, 3215, 3187, 3187, 3187, 3187, 3187, 3187, 3187, 3187, 3187, 3187, 3187, 3187, 3152, 3152, 3152, 3152, 3152, 3152, 3152, 3152, 3152, 3152, 3152, 3152, 3152, 3125, 3125, 3125, 3125, 3125, 3125, 3125, 3125, 3125, 3125, 3125, 3125, 3125, 3090, 3090, 3090, 3090, 3090, 3090, 3090, 3090, 3090, 3090, 3090, 3090, 3090, 3062, 3062, 3062, 3062, 3062, 3062, 3062, 3062, 3062, 3062, 3062, 3062, 3062, 3062, 3027, 3027, 3027, 3027, 3027, 3027, 3027, 3027, 3027, 3027, 3027, 3027, 3027, 2999, 2999, 2999, 2999, 2999, 2999, 2999, 2999, 2999, 2999, 2999, 2999, 2999, 2964, 2964, 2964, 2964, 2964, 2964, 2964, 2964, 2964, 2964, 2964, 2964, 2964, 2937, 2937, 2937, 2937, 2937, 2937, 2937, 2937, 2937, 2937, 2937, 2937, 2937, 2937, 2902, 2902, 2902, 2902, 2902, 2902, 2902, 2902, 2902, 2902, 2902, 2902, 2902, 2874, 2874, 2874, 2874, 2874, 2874, 2874, 2874, 2874, 2874, 2874, 2874, 2874, 2874, 2846, 2846, 2846, 2846, 2846, 2846, 2846, 2846, 2846, 2846, 2846, 2846, 2846, 2846, 2811, 2811, 2811, 2811, 2811, 2811, 2811, 2811, 2811, 2811, 2811, 2811, 2811, 2783, 2783, 2783, 2783, 2783, 2783, 2783, 2783, 2783, 2783, 2783, 2783, 2783, 2783, 2748, 2748, 2748, 2748, 2748, 2748, 2748, 2748, 2748, 2748, 2748, 2748, 2748, 2748, 2720, 2720, 2720, 2720, 2720, 2720, 2720, 2720, 2720, 2720, 2720, 2720, 2720, 2720, 2685, 2685, 2685, 2685, 2685, 2685, 2685, 2685, 2685, 2685, 2685, 2685, 2685, 2685, 2657, 2657, 2657, 2657, 2657, 2657, 2657, 2657, 2657, 2657, 2657, 2657, 2657, 2657, 2622, 2622, 2622, 2622, 2622, 2622, 2622, 2622, 2622, 2622, 2622, 2622, 2622, 2622, 2594, 2594, 2594, 2594, 2594, 2594, 2594, 2594, 2594, 2594, 2594, 2594, 2594, 2594, 2594, 2559, 2559, 2559, 2559, 2559, 2559, 2559, 2559, 2559, 2559, 2559, 2559, 2559, 2559, 2531, 2531, 2531, 2531, 2531, 2531, 2531, 2531, 2531, 2531, 2531, 2531, 2531, 2531, 2496, 2496, 2496, 2496, 2496, 2496, 2496, 2496, 2496, 2496, 2496, 2496, 2496, 2496, 2496, 2468, 2468, 2468, 2468, 2468, 2468, 2468, 2468, 2468, 2468, 2468, 2468, 2468, 2468, 2468, 2433, 2433, 2433, 2433, 2433, 2433, 2433, 2433, 2433, 2433, 2433, 2433, 2433, 2433, 2405, 2405, 2405, 2405, 2405, 2405, 2405, 2405, 2405, 2405, 2405, 2405, 2405, 2405, 2405, 2370, 2370, 2370, 2370, 2370, 2370, 2370, 2370, 2370, 2370, 2370, 2370, 2370, 2370, 2370, 2342, 2342, 2342, 2342, 2342, 2342, 2342, 2342, 2342, 2342, 2342, 2342, 2342, 2342, 2342, 2307, 2307, 2307, 2307, 2307, 2307, 2307, 2307, 2307, 2307, 2307, 2307, 2307, 2307, 2307, 2278, 2278, 2278, 2278, 2278, 2278, 2278, 2278, 2278, 2278, 2278, 2278, 2278, 2278, 2278, 2278, 2243, 2243, 2243, 2243, 2243, 2243, 2243, 2243, 2243, 2243, 2243, 2243, 2243, 2243, 2243, 2215, 2215, 2215, 2215, 2215, 2215, 2215, 2215, 2215, 2215, 2215, 2215, 2215, 2215, 2215, 2180, 2180, 2180, 2180, 2180, 2180, 2180, 2180, 2180, 2180, 2180, 2180, 2180, 2180, 2180, 2180, 2152, 2152, 2152, 2152, 2152, 2152, 2152, 2152, 2152, 2152, 2152, 2152, 2152, 2152, 2152, 2152, 2116, 2116, 2116, 2116, 2116, 2116, 2116, 2116, 2116, 2116, 2116, 2116, 2116, 2116, 2116, 2088, 2088, 2088, 2088, 2088, 2088, 2088, 2088, 2088, 2088, 2088, 2088, 2088, 2088, 2088, 2088, 2053, 2053, 2053, 2053, 2053, 2053, 2053, 2053, 2053, 2053, 2053, 2053, 2053, 2053, 2053, 2053, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 1989, 1989, 1989, 1989, 1989, 1989, 1989, 1989, 1989, 1989, 1989, 1989, 1989, 1989, 1989, 1989, 1961, 1961, 1961, 1961, 1961, 1961, 1961, 1961, 1961, 1961, 1961, 1961, 1961, 1961, 1961, 1961, 1926, 1926, 1926, 1926, 1926, 1926, 1926, 1926, 1926, 1926, 1926, 1926, 1926, 1926, 1926, 1926, 1926, 1898, 1898, 1898, 1898, 1898, 1898, 1898, 1898, 1898, 1898, 1898, 1898, 1898, 1898, 1898, 1898, 1898, 1862, 1862, 1862, 1862, 1862, 1862, 1862, 1862, 1862, 1862, 1862, 1862, 1862, 1862, 1862, 1862, 1862, 1834, 1834, 1834, 1834, 1834, 1834, 1834, 1834, 1834, 1834, 1834, 1834, 1834, 1834, 1834, 1834, 1834, 1799, 1799, 1799, 1799, 1799, 1799, 1799, 1799, 1799, 1799, 1799, 1799, 1799, 1799, 1799, 1799, 1799, 1770, 1770, 1770, 1770, 1770, 1770, 1770, 1770, 1770, 1770, 1770, 1770, 1770, 1770, 1770, 1770, 1770, 1735, 1735, 1735, 1735, 1735, 1735, 1735, 1735, 1735, 1735, 1735, 1735, 1735, 1735, 1735, 1735, 1735, 1735, 1707, 1707, 1707, 1707, 1707, 1707, 1707, 1707, 1707, 1707, 1707, 1707, 1707, 1707, 1707, 1707, 1707, 1671, 1671, 1671, 1671, 1671, 1671, 1671, 1671, 1671, 1671, 1671, 1671, 1671, 1671, 1671, 1671, 1671, 1671, 1643, 1643, 1643, 1643, 1643, 1643, 1643, 1643, 1643, 1643, 1643, 1643, 1643, 1643, 1643, 1643, 1643, 1643, 1607, 1607, 1607, 1607, 1607, 1607, 1607, 1607, 1607, 1607, 1607, 1607, 1607, 1607, 1607, 1607, 1607, 1607, 1579, 1579, 1579, 1579, 1579, 1579, 1579, 1579, 1579, 1579, 1579, 1579, 1579, 1579, 1579, 1579, 1579, 1579, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1543, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1515, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1479, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1451, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1422, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1387, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1358, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1323, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1294, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1259, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1230, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1194, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1166, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1130, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1102, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1066, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1037, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 937, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 908, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 873, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 844, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 808, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 779, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 743, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 715, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 679, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 650, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 614, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 585, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 549, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 484, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 456, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 420, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 391, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 326, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 261, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 225, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 72000, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71971, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71935, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71906, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71870, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71841, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71804, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71775, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71739, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71710, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71674, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71645, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71609, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71580, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71544, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71516, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71480, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71451, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71415, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71386, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71350, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71321, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71285, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71257, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71221, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71192, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71156, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71127, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71092, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71063, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 71027, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70998, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70963, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70934, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70898, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70870, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70834, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70806, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70770, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70741, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70706, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70677, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70642, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70613, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70578, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70549, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70521, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70485, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70457, 70421, 70421, 70421, 70421, 70421, 70421, 70421, 70421, 70421, 70421, 70421, 70421, 70421, 70421, 70421, 70421, 70421, 70421, 70393, 70393, 70393, 70393, 70393, 70393, 70393, 70393, 70393, 70393, 70393, 70393, 70393, 70393, 70393, 70393, 70393, 70393, 70357, 70357, 70357, 70357, 70357, 70357, 70357, 70357, 70357, 70357, 70357, 70357, 70357, 70357, 70357, 70357, 70357, 70357, 70329, 70329, 70329, 70329, 70329, 70329, 70329, 70329, 70329, 70329, 70329, 70329, 70329, 70329, 70329, 70329, 70329, 70329, 70293, 70293, 70293, 70293, 70293, 70293, 70293, 70293, 70293, 70293, 70293, 70293, 70293, 70293, 70293, 70293, 70293, 70265, 70265, 70265, 70265, 70265, 70265, 70265, 70265, 70265, 70265, 70265, 70265, 70265, 70265, 70265, 70265, 70265, 70265, 70230, 70230, 70230, 70230, 70230, 70230, 70230, 70230, 70230, 70230, 70230, 70230, 70230, 70230, 70230, 70230, 70230, 70201, 70201, 70201, 70201, 70201, 70201, 70201, 70201, 70201, 70201, 70201, 70201, 70201, 70201, 70201, 70201, 70201, 70166, 70166, 70166, 70166, 70166, 70166, 70166, 70166, 70166, 70166, 70166, 70166, 70166, 70166, 70166, 70166, 70166, 70138, 70138, 70138, 70138, 70138, 70138, 70138, 70138, 70138, 70138, 70138, 70138, 70138, 70138, 70138, 70138, 70138, 70102, 70102, 70102, 70102, 70102, 70102, 70102, 70102, 70102, 70102, 70102, 70102, 70102, 70102, 70102, 70102, 70102, 70074, 70074, 70074, 70074, 70074, 70074, 70074, 70074, 70074, 70074, 70074, 70074, 70074, 70074, 70074, 70074, 70074, 70039, 70039, 70039, 70039, 70039, 70039, 70039, 70039, 70039, 70039, 70039, 70039, 70039, 70039, 70039, 70039, 70011, 70011, 70011, 70011, 70011, 70011, 70011, 70011, 70011, 70011, 70011, 70011, 70011, 70011, 70011, 70011, 69975, 69975, 69975, 69975, 69975, 69975, 69975, 69975, 69975, 69975, 69975, 69975, 69975, 69975, 69975, 69975, 69975, 69947, 69947, 69947, 69947, 69947, 69947, 69947, 69947, 69947, 69947, 69947, 69947, 69947, 69947, 69947, 69947, 69912, 69912, 69912, 69912, 69912, 69912, 69912, 69912, 69912, 69912, 69912, 69912, 69912, 69912, 69912, 69912, 69884, 69884, 69884, 69884, 69884, 69884, 69884, 69884, 69884, 69884, 69884, 69884, 69884, 69884, 69884, 69848, 69848, 69848, 69848, 69848, 69848, 69848, 69848, 69848, 69848, 69848, 69848, 69848, 69848, 69848, 69848, 69820, 69820, 69820, 69820, 69820, 69820, 69820, 69820, 69820, 69820, 69820, 69820, 69820, 69820, 69820, 69820, 69785, 69785, 69785, 69785, 69785, 69785, 69785, 69785, 69785, 69785, 69785, 69785, 69785, 69785, 69785, 69757, 69757, 69757, 69757, 69757, 69757, 69757, 69757, 69757, 69757, 69757, 69757, 69757, 69757, 69757, 69722, 69722, 69722, 69722, 69722, 69722, 69722, 69722, 69722, 69722, 69722, 69722, 69722, 69722, 69722, 69722, 69693, 69693, 69693, 69693, 69693, 69693, 69693, 69693, 69693, 69693, 69693, 69693, 69693, 69693, 69693, 69658, 69658, 69658, 69658, 69658, 69658, 69658, 69658, 69658, 69658, 69658, 69658, 69658, 69658, 69658, 69630, 69630, 69630, 69630, 69630, 69630, 69630, 69630, 69630, 69630, 69630, 69630, 69630, 69630, 69630, 69595, 69595, 69595, 69595, 69595, 69595, 69595, 69595, 69595, 69595, 69595, 69595, 69595, 69595, 69595, 69567, 69567, 69567, 69567, 69567, 69567, 69567, 69567, 69567, 69567, 69567, 69567, 69567, 69567, 69532, 69532, 69532, 69532, 69532, 69532, 69532, 69532, 69532, 69532, 69532, 69532, 69532, 69532, 69532, 69504, 69504, 69504, 69504, 69504, 69504, 69504, 69504, 69504, 69504, 69504, 69504, 69504, 69504, 69504, 69469, 69469, 69469, 69469, 69469, 69469, 69469, 69469, 69469, 69469, 69469, 69469, 69469, 69469, 69441, 69441, 69441, 69441, 69441, 69441, 69441, 69441, 69441, 69441, 69441, 69441, 69441, 69441, 69406, 69406, 69406, 69406, 69406, 69406, 69406, 69406, 69406, 69406, 69406, 69406, 69406, 69406, 69406, 69378, 69378, 69378, 69378, 69378, 69378, 69378, 69378, 69378, 69378, 69378, 69378, 69378, 69378, 69343, 69343, 69343, 69343, 69343, 69343, 69343, 69343, 69343, 69343, 69343, 69343, 69343, 69343, 69315, 69315, 69315, 69315, 69315, 69315, 69315, 69315, 69315, 69315, 69315, 69315, 69315, 69315, 69280, 69280, 69280, 69280, 69280, 69280, 69280, 69280, 69280, 69280, 69280, 69280, 69280, 69280, 69252, 69252, 69252, 69252, 69252, 69252, 69252, 69252, 69252, 69252, 69252, 69252, 69252, 69252, 69217, 69217, 69217, 69217, 69217, 69217, 69217, 69217, 69217, 69217, 69217, 69217, 69217, 69217, 69189, 69189, 69189, 69189, 69189, 69189, 69189, 69189, 69189, 69189, 69189, 69189, 69189, 69154, 69154, 69154, 69154, 69154, 69154, 69154, 69154, 69154, 69154, 69154, 69154, 69154, 69154, 69126, 69126, 69126, 69126, 69126, 69126, 69126, 69126, 69126, 69126, 69126, 69126, 69126, 69126, 69098, 69098, 69098, 69098, 69098, 69098, 69098, 69098, 69098, 69098, 69098, 69098, 69098, 69063, 69063, 69063, 69063, 69063, 69063, 69063, 69063, 69063, 69063, 69063, 69063, 69063, 69063, 69036, 69036, 69036, 69036, 69036, 69036, 69036, 69036, 69036, 69036, 69036, 69036, 69036, 69001, 69001, 69001, 69001, 69001, 69001, 69001, 69001, 69001, 69001, 69001, 69001, 69001, 68973, 68973, 68973, 68973, 68973, 68973, 68973, 68973, 68973, 68973, 68973, 68973, 68973, 68938, 68938, 68938, 68938, 68938, 68938, 68938, 68938, 68938, 68938, 68938, 68938, 68938, 68938, 68910, 68910, 68910, 68910, 68910, 68910, 68910, 68910, 68910, 68910, 68910, 68910, 68910, 68875, 68875, 68875, 68875, 68875, 68875, 68875, 68875, 68875, 68875, 68875, 68875, 68875, 68848, 68848, 68848, 68848, 68848, 68848, 68848, 68848, 68848, 68848, 68848, 68848, 68848, 68813, 68813, 68813, 68813, 68813, 68813, 68813, 68813, 68813, 68813, 68813, 68813, 68785, 68785, 68785, 68785, 68785, 68785, 68785, 68785, 68785, 68785, 68785, 68785, 68785, 68750, 68750, 68750, 68750, 68750, 68750, 68750, 68750, 68750, 68750, 68750, 68750, 68750, 68723, 68723, 68723, 68723, 68723, 68723, 68723, 68723, 68723, 68723, 68723, 68723, 68723, 68688, 68688, 68688, 68688, 68688, 68688, 68688, 68688, 68688, 68688, 68688, 68688, 68660, 68660, 68660, 68660, 68660, 68660, 68660, 68660, 68660, 68660, 68660, 68660, 68660, 68626, 68626, 68626, 68626, 68626, 68626, 68626, 68626, 68626, 68626, 68626, 68626, 68598, 68598, 68598, 68598, 68598, 68598, 68598, 68598, 68598, 68598, 68598, 68598, 68598, 68563, 68563, 68563, 68563, 68563, 68563, 68563, 68563, 68563, 68563, 68563, 68563, 68535, 68535, 68535, 68535, 68535, 68535, 68535, 68535, 68535, 68535, 68535, 68535, 68535, 68501, 68501, 68501, 68501, 68501, 68501, 68501, 68501, 68501, 68501, 68501, 68501, 68473, 68473, 68473, 68473, 68473, 68473, 68473, 68473, 68473, 68473, 68473, 68473, 68439, 68439, 68439, 68439, 68439, 68439, 68439, 68439, 68439, 68439, 68439, 68439, 68411, 68411, 68411, 68411, 68411, 68411, 68411, 68411, 68411, 68411, 68411, 68411, 68376, 68376, 68376, 68376, 68376, 68376, 68376, 68376, 68376, 68376, 68376, 68376, 68349, 68349, 68349, 68349, 68349, 68349, 68349, 68349, 68349, 68349, 68349, 68349, 68314, 68314, 68314, 68314, 68314, 68314, 68314, 68314, 68314, 68314, 68314, 68314, 68287, 68287, 68287, 68287, 68287, 68287, 68287, 68287, 68287, 68287, 68287, 68287, 68252, 68252, 68252, 68252, 68252, 68252, 68252, 68252, 68252, 68252, 68252, 68252, 68225, 68225, 68225, 68225, 68225, 68225, 68225, 68225, 68225, 68225, 68225, 68225, 68190, 68190, 68190, 68190, 68190, 68190, 68190, 68190, 68190, 68190, 68190, 68190, 68163, 68163, 68163, 68163, 68163, 68163, 68163, 68163, 68163, 68163, 68163, 68163, 68128, 68128, 68128, 68128, 68128, 68128, 68128, 68128, 68128, 68128, 68128, 68101, 68101, 68101, 68101, 68101, 68101, 68101, 68101, 68101, 68101, 68101, 68101, 68066, 68066, 68066, 68066, 68066, 68066, 68066, 68066, 68066, 68066, 68066, 68039, 68039, 68039, 68039, 68039, 68039, 68039, 68039, 68039, 68039, 68039, 68039, 68004, 68004, 68004, 68004, 68004, 68004, 68004, 68004, 68004, 68004, 68004, 67977, 67977, 67977, 67977, 67977, 67977, 67977, 67977, 67977, 67977, 67977, 67977, 67942, 67942, 67942, 67942, 67942, 67942, 67942, 67942, 67942, 67942, 67942, 67915, 67915, 67915, 67915, 67915, 67915, 67915, 67915, 67915, 67915, 67915, 67915, 67881, 67881, 67881, 67881, 67881, 67881, 67881, 67881, 67881, 67881, 67881, 67853, 67853, 67853, 67853, 67853, 67853, 67853, 67853, 67853, 67853, 67853, 67819, 67819, 67819, 67819, 67819, 67819, 67819, 67819, 67819, 67819, 67819, 67791, 67791, 67791, 67791, 67791, 67791, 67791, 67791, 67791, 67791, 67791, 67791, 67764, 67764, 67764, 67764, 67764, 67764, 67764, 67764, 67764, 67764, 67764, 67730, 67730, 67730, 67730, 67730, 67730, 67730, 67730, 67730, 67730, 67730, 67702, 67702, 67702, 67702, 67702, 67702, 67702, 67702, 67702, 67702, 67702, 67668, 67668, 67668, 67668, 67668, 67668, 67668, 67668, 67668, 67668, 67668, 67641, 67641, 67641, 67641, 67641, 67641, 67641, 67641, 67641, 67641, 67641, 67607, 67607, 67607, 67607, 67607, 67607, 67607, 67607, 67607, 67607, 67607, 67579, 67579, 67579, 67579, 67579, 67579, 67579, 67579, 67579, 67579, 67579, 67545, 67545, 67545, 67545, 67545, 67545, 67545, 67545, 67545, 67545, 67545, 67518, 67518, 67518, 67518, 67518, 67518, 67518, 67518, 67518, 67518, 67518, 67484, 67484, 67484, 67484, 67484, 67484, 67484, 67484, 67484, 67484, 67456, 67456, 67456, 67456, 67456, 67456, 67456, 67456, 67456, 67456, 67456, 67422, 67422, 67422, 67422, 67422, 67422, 67422, 67422, 67422, 67422, 67422, 67395, 67395, 67395, 67395, 67395, 67395, 67395, 67395, 67395, 67395, 67395, 67361, 67361, 67361, 67361, 67361, 67361, 67361, 67361, 67361, 67361, 67333, 67333, 67333, 67333, 67333, 67333, 67333, 67333, 67333, 67333, 67333, 67299, 67299, 67299, 67299, 67299, 67299, 67299, 67299, 67299, 67299, 67272, 67272, 67272, 67272, 67272, 67272, 67272, 67272, 67272, 67272, 67272, 67238, 67238, 67238, 67238, 67238, 67238, 67238, 67238, 67238, 67238, 67211, 67211, 67211, 67211, 67211, 67211, 67211, 67211, 67211, 67211, 67211, 67177, 67177, 67177, 67177, 67177, 67177, 67177, 67177, 67177, 67177, 67150, 67150, 67150, 67150, 67150, 67150, 67150, 67150, 67150, 67150, 67150, 67116, 67116, 67116, 67116, 67116, 67116, 67116, 67116, 67116, 67116, 67088, 67088, 67088, 67088, 67088, 67088, 67088, 67088, 67088, 67088, 67055, 67055, 67055, 67055, 67055, 67055, 67055, 67055, 67055, 67055, 67055, 67027, 67027, 67027, 67027, 67027, 67027, 67027, 67027, 67027, 67027, 66993, 66993, 66993, 66993, 66993, 66993, 66993, 66993, 66993, 66993, 66966, 66966, 66966, 66966, 66966, 66966, 66966, 66966, 66966, 66966, 66966, 66932, 66932, 66932, 66932, 66932, 66932, 66932, 66932, 66932, 66932, 66905, 66905, 66905, 66905, 66905, 66905, 66905, 66905, 66905, 66905, 66871, 66871, 66871, 66871, 66871, 66871, 66871, 66871, 66871, 66871, 66844, 66844, 66844, 66844, 66844, 66844, 66844, 66844, 66844, 66844, 66810, 66810, 66810, 66810, 66810, 66810, 66810, 66810, 66810, 66810, 66783, 66783, 66783, 66783, 66783, 66783, 66783, 66783, 66783, 66783, 66750, 66750, 66750, 66750, 66750, 66750, 66750, 66750, 66750, 66750, 66722, 66722, 66722, 66722, 66722, 66722, 66722, 66722, 66722, 66722, 66689, 66689, 66689, 66689, 66689, 66689, 66689, 66689, 66689, 66689, 66662, 66662, 66662, 66662, 66662, 66662, 66662, 66662, 66662, 66662, 66628, 66628, 66628, 66628, 66628, 66628, 66628, 66628, 66628, 66628, 66601, 66601, 66601, 66601, 66601, 66601, 66601, 66601, 66601, 66601, 66567, 66567, 66567, 66567, 66567, 66567, 66567, 66567, 66567, 66567, 66540, 66540, 66540, 66540, 66540, 66540, 66540, 66540, 66540, 66506, 66506, 66506, 66506, 66506, 66506, 66506, 66506, 66506, 66506, 66479, 66479, 66479, 66479, 66479, 66479, 66479, 66479, 66479, 66479, 66446, 66446, 66446, 66446, 66446, 66446, 66446, 66446, 66446, 66446, 66419, 66419, 66419, 66419, 66419, 66419, 66419, 66419, 66419, 66392, 66392, 66392, 66392, 66392, 66392, 66392, 66392, 66392, 66392, 66358, 66358, 66358, 66358, 66358, 66358, 66358, 66358, 66358, 66358, 66331, 66331, 66331, 66331, 66331, 66331, 66331, 66331, 66331, 66298, 66298, 66298, 66298, 66298, 66298, 66298, 66298, 66298, 66298, 66271, 66271, 66271, 66271, 66271, 66271, 66271, 66271, 66271, 66271, 66237, 66237, 66237, 66237, 66237, 66237, 66237, 66237, 66237, 66210, 66210, 66210, 66210, 66210, 66210, 66210, 66210, 66210, 66210, 66177, 66177, 66177, 66177, 66177, 66177, 66177, 66177, 66177, 66150, 66150, 66150, 66150, 66150, 66150, 66150, 66150, 66150, 66150, 66116, 66116, 66116, 66116, 66116, 66116, 66116, 66116, 66116, 66089, 66089, 66089, 66089, 66089, 66089, 66089, 66089, 66089, 66056, 66056, 66056, 66056, 66056, 66056, 66056, 66056, 66056, 66056, 66029, 66029, 66029, 66029, 66029, 66029, 66029, 66029, 66029, 65995, 65995, 65995, 65995, 65995, 65995, 65995, 65995, 65995, 65995, 65969, 65969, 65969, 65969, 65969, 65969, 65969, 65969, 65969, 65935, 65935, 65935, 65935, 65935, 65935, 65935, 65935, 65935, 65908, 65908, 65908, 65908, 65908, 65908, 65908, 65908, 65908, 65875, 65875, 65875, 65875, 65875, 65875, 65875, 65875, 65875, 65875, 65848, 65848, 65848, 65848, 65848, 65848, 65848, 65848, 65848, 65815, 65815, 65815, 65815, 65815, 65815, 65815, 65815, 65815, 65788, 65788, 65788, 65788, 65788, 65788, 65788, 65788, 65788, 65755, 65755, 65755, 65755, 65755, 65755, 65755, 65755, 65755, 65728, 65728, 65728, 65728, 65728, 65728, 65728, 65728, 65728, 65728, 65695, 65695, 65695, 65695, 65695, 65695, 65695, 65695, 65695, 65668, 65668, 65668, 65668, 65668, 65668, 65668, 65668, 65668, 65634, 65634, 65634, 65634, 65634, 65634, 65634, 65634, 65634, 65608, 65608, 65608, 65608, 65608, 65608, 65608, 65608, 65608, 65574, 65574, 65574, 65574, 65574, 65574, 65574, 65574, 65574, 65548, 65548, 65548, 65548, 65548, 65548, 65548, 65548, 65548, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65455, 65455, 65455, 65455, 65455, 65455, 65455, 65455, 65455, 65428, 65428, 65428, 65428, 65428, 65428, 65428, 65428, 65428, 65395, 65395, 65395, 65395, 65395, 65395, 65395, 65395, 65395, 65368, 65368, 65368, 65368, 65368, 65368, 65368, 65368, 65368, 65335, 65335, 65335, 65335, 65335, 65335, 65335, 65335, 65308, 65308, 65308, 65308, 65308, 65308, 65308, 65308, 65308, 65275, 65275, 65275, 65275, 65275, 65275, 65275, 65275, 65275, 65248, 65248, 65248, 65248, 65248, 65248, 65248, 65248, 65248, 65215, 65215, 65215, 65215, 65215, 65215, 65215, 65215, 65215, 65189, 65189, 65189, 65189, 65189, 65189, 65189, 65189, 65189, 65156, 65156, 65156, 65156, 65156, 65156, 65156, 65156, 65129, 65129, 65129, 65129, 65129, 65129, 65129, 65129, 65129, 65096, 65096, 65096, 65096, 65096, 65096, 65096, 65096, 65096, 65069, 65069, 65069, 65069, 65069, 65069, 65069, 65069, 65043, 65043, 65043, 65043, 65043, 65043, 65043, 65043, 65043, 65010, 65010, 65010, 65010, 65010, 65010, 65010, 65010, 65010, 64983, 64983, 64983, 64983, 64983, 64983, 64983, 64983, 64950, 64950, 64950, 64950, 64950, 64950, 64950, 64950, 64950, 64924, 64924, 64924, 64924, 64924, 64924, 64924, 64924, 64924, 64891, 64891, 64891, 64891, 64891, 64891, 64891, 64891, 64864, 64864, 64864, 64864, 64864, 64864, 64864, 64864, 64864, 64831, 64831, 64831, 64831, 64831, 64831, 64831, 64831, 64805, 64805, 64805, 64805, 64805, 64805, 64805, 64805, 64805, 64772, 64772, 64772, 64772, 64772, 64772, 64772, 64772, 64746, 64746, 64746, 64746, 64746, 64746, 64746, 64746, 64746, 64713, 64713, 64713, 64713, 64713, 64713, 64713, 64713, 64686, 64686, 64686, 64686, 64686, 64686, 64686, 64686, 64686, 64653, 64653, 64653, 64653, 64653, 64653, 64653, 64653, 64627, 64627, 64627, 64627, 64627, 64627, 64627, 64627, 64627, 64594, 64594, 64594, 64594, 64594, 64594, 64594, 64594, 64568, 64568, 64568, 64568, 64568, 64568, 64568, 64568, 64535, 64535, 64535, 64535, 64535, 64535, 64535, 64535, 64535, 64508, 64508, 64508, 64508, 64508, 64508, 64508, 64508, 64475, 64475, 64475, 64475, 64475, 64475, 64475, 64475, 64449, 64449, 64449, 64449, 64449, 64449, 64449, 64449, 64449, 64416, 64416, 64416, 64416, 64416, 64416, 64416, 64416, 64390, 64390, 64390, 64390, 64390, 64390, 64390, 64390, 64357, 64357, 64357, 64357, 64357, 64357, 64357, 64357, 64357, 64331, 64331, 64331, 64331, 64331, 64331, 64331, 64331, 64298, 64298, 64298, 64298, 64298, 64298, 64298, 64298, 64272, 64272, 64272, 64272, 64272, 64272, 64272, 64272, 64239, 64239, 64239, 64239, 64239, 64239, 64239, 64239, 64239, 64213, 64213, 64213, 64213, 64213, 64213, 64213, 64213, 64180, 64180, 64180, 64180, 64180, 64180, 64180, 64180, 64154, 64154, 64154, 64154, 64154, 64154, 64154, 64154, 64121, 64121, 64121, 64121, 64121, 64121, 64121, 64121, 64095, 64095, 64095, 64095, 64095, 64095, 64095, 64095, 64062, 64062, 64062, 64062, 64062, 64062, 64062, 64062, 64036, 64036, 64036, 64036, 64036, 64036, 64036, 64036, 64036, 64003, 64003, 64003, 64003, 64003, 64003, 64003, 64003, 63977, 63977, 63977, 63977, 63977, 63977, 63977, 63977, 63944, 63944, 63944, 63944, 63944, 63944, 63944, 63944, 63918, 63918, 63918, 63918, 63918, 63918, 63918, 63918, 63886, 63886, 63886, 63886, 63886, 63886, 63886, 63886, 63860, 63860, 63860, 63860, 63860, 63860, 63860, 63860, 63827, 63827, 63827, 63827, 63827, 63827, 63827, 63827, 63801, 63801, 63801, 63801, 63801, 63801, 63801, 63801, 63768, 63768, 63768, 63768, 63768, 63768, 63768, 63768, 63742, 63742, 63742, 63742, 63742, 63742, 63742, 63742, 63716, 63716, 63716, 63716, 63716, 63716, 63716, 63716, 63684, 63684, 63684, 63684, 63684, 63684, 63684, 63684, 63657, 63657, 63657, 63657, 63657, 63657, 63657, 63625, 63625, 63625, 63625, 63625, 63625, 63625, 63625, 63599, 63599, 63599, 63599, 63599, 63599, 63599, 63599, 63566, 63566, 63566, 63566, 63566, 63566, 63566, 63566, 63540, 63540, 63540, 63540, 63540, 63540, 63540, 63540, 63508, 63508, 63508, 63508, 63508, 63508, 63508, 63508, 63482, 63482, 63482, 63482, 63482, 63482, 63482, 63482, 63449, 63449, 63449, 63449, 63449, 63449, 63449, 63423, 63423, 63423, 63423, 63423, 63423, 63423, 63423, 63391, 63391, 63391, 63391, 63391, 63391, 63391, 63391, 63365, 63365, 63365, 63365, 63365, 63365, 63365, 63365, 63332, 63332, 63332, 63332, 63332, 63332, 63332, 63332, 63307, 63307, 63307, 63307, 63307, 63307, 63307, 63274, 63274, 63274, 63274, 63274, 63274, 63274, 63274, 63248, 63248, 63248, 63248, 63248, 63248, 63248, 63248, 63216, 63216, 63216, 63216, 63216, 63216, 63216, 63190, 63190, 63190, 63190, 63190, 63190, 63190, 63190, 63158, 63158, 63158, 63158, 63158, 63158, 63158, 63158, 63132, 63132, 63132, 63132, 63132, 63132, 63132, 63099, 63099, 63099, 63099, 63099, 63099, 63099, 63099, 63073, 63073, 63073, 63073, 63073, 63073, 63073, 63073, 63041, 63041, 63041, 63041, 63041, 63041, 63041, 63015, 63015, 63015, 63015, 63015, 63015, 63015, 63015, 62983, 62983, 62983, 62983, 62983, 62983, 62983, 62983, 62957, 62957, 62957, 62957, 62957, 62957, 62957, 62925, 62925, 62925, 62925, 62925, 62925, 62925, 62925, 62899, 62899, 62899, 62899, 62899, 62899, 62899, 62867, 62867, 62867, 62867, 62867, 62867, 62867, 62867, 62841, 62841, 62841, 62841, 62841, 62841, 62841, 62809, 62809, 62809, 62809, 62809, 62809, 62809, 62809, 62783, 62783, 62783, 62783, 62783, 62783, 62783, 62751, 62751, 62751, 62751, 62751, 62751, 62751, 62751, 62725, 62725, 62725, 62725, 62725, 62725, 62725, 62693, 62693, 62693, 62693, 62693, 62693, 62693, 62693, 62667, 62667, 62667, 62667, 62667, 62667, 62667, 62635, 62635, 62635, 62635, 62635, 62635, 62635, 62635, 62609, 62609, 62609, 62609, 62609, 62609, 62609, 62577, 62577, 62577, 62577, 62577, 62577, 62577, 62577, 62551, 62551, 62551, 62551, 62551, 62551, 62551, 62519, 62519, 62519, 62519, 62519, 62519, 62519, 62519, 62493, 62493, 62493, 62493, 62493, 62493, 62493, 62468, 62468, 62468, 62468, 62468, 62468, 62468, 62436, 62436, 62436, 62436, 62436, 62436, 62436, 62436, 62410, 62410, 62410, 62410, 62410, 62410, 62410, 62378, 62378, 62378, 62378, 62378, 62378, 62378, 62352, 62352, 62352, 62352, 62352, 62352, 62352, 62352, 62320, 62320, 62320, 62320, 62320, 62320, 62320, 62294, 62294, 62294, 62294, 62294, 62294, 62294, 62262, 62262, 62262, 62262, 62262, 62262, 62262, 62262, 62237, 62237, 62237, 62237, 62237, 62237, 62237, 62205, 62205, 62205, 62205, 62205, 62205, 62205, 62179, 62179, 62179, 62179, 62179, 62179, 62179, 62179, 62147, 62147, 62147, 62147, 62147, 62147, 62147, 62122, 62122, 62122, 62122, 62122, 62122, 62122, 62090, 62090, 62090, 62090, 62090, 62090, 62090, 62064, 62064, 62064, 62064, 62064, 62064, 62064, 62064, 62032, 62032, 62032, 62032, 62032, 62032, 62032, 62006, 62006, 62006, 62006, 62006, 62006, 62006, 61975, 61975, 61975, 61975, 61975, 61975, 61975, 61949, 61949, 61949, 61949, 61949, 61949, 61949, 61949, 61917, 61917, 61917, 61917, 61917, 61917, 61917, 61892, 61892, 61892, 61892, 61892, 61892, 61892, 61860, 61860, 61860, 61860, 61860, 61860, 61860, 61834, 61834, 61834, 61834, 61834, 61834, 61834, 61802, 61802, 61802, 61802, 61802, 61802, 61802, 61777, 61777, 61777, 61777, 61777, 61777, 61777, 61745, 61745, 61745, 61745, 61745, 61745, 61745, 61745, 61719, 61719, 61719, 61719, 61719, 61719, 61719, 61688, 61688, 61688, 61688, 61688, 61688, 61688, 61662, 61662, 61662, 61662, 61662, 61662, 61662, 61630, 61630, 61630, 61630, 61630, 61630, 61630, 61605, 61605, 61605, 61605, 61605, 61605, 61605, 61573, 61573, 61573, 61573, 61573, 61573, 61573, 61548, 61548, 61548, 61548, 61548, 61548, 61548, 61516, 61516, 61516, 61516, 61516, 61516, 61516, 61491, 61491, 61491, 61491, 61491, 61491, 61491, 61459, 61459, 61459, 61459, 61459, 61459, 61459, 61433, 61433, 61433, 61433, 61433, 61433, 61433, 61402, 61402, 61402, 61402, 61402, 61402, 61402, 61376, 61376, 61376, 61376, 61376, 61376, 61376, 61345, 61345, 61345, 61345, 61345, 61345, 61345, 61319, 61319, 61319, 61319, 61319, 61319, 61319, 61288, 61288, 61288, 61288, 61288, 61288, 61288, 61262, 61262, 61262, 61262, 61262, 61262, 61262, 61231, 61231, 61231, 61231, 61231, 61231, 61231, 61205, 61205, 61205, 61205, 61205, 61205, 61205, 61180, 61180, 61180, 61180, 61180, 61180, 61180, 61148, 61148, 61148, 61148, 61148, 61148, 61148, 61123, 61123, 61123, 61123, 61123, 61123, 61123, 61091, 61091, 61091, 61091, 61091, 61091, 61091, 61066, 61066, 61066, 61066, 61066, 61066, 61066, 61034, 61034, 61034, 61034, 61034, 61034, 61009, 61009, 61009, 61009, 61009, 61009, 61009, 60978, 60978, 60978, 60978, 60978, 60978, 60978, 60952, 60952, 60952, 60952, 60952, 60952, 60952, 60921, 60921, 60921, 60921, 60921, 60921, 60921, 60896, 60896, 60896, 60896, 60896, 60896, 60896, 60864, 60864, 60864, 60864, 60864, 60864, 60864, 60839, 60839, 60839, 60839, 60839, 60839, 60807, 60807, 60807, 60807, 60807, 60807, 60807, 60782, 60782, 60782, 60782, 60782, 60782, 60782, 60751, 60751, 60751, 60751, 60751, 60751, 60751, 60725, 60725, 60725, 60725, 60725, 60725, 60725, 60694, 60694, 60694, 60694, 60694, 60694, 60669, 60669, 60669, 60669, 60669, 60669, 60669, 60637, 60637, 60637, 60637, 60637, 60637, 60637, 60612, 60612, 60612, 60612, 60612, 60612, 60612, 60581, 60581, 60581, 60581, 60581, 60581, 60556, 60556, 60556, 60556, 60556, 60556, 60556, 60524, 60524, 60524, 60524, 60524, 60524, 60524, 60499, 60499, 60499, 60499, 60499, 60499, 60499, 60468, 60468, 60468, 60468, 60468, 60468, 60442, 60442, 60442, 60442, 60442, 60442, 60442, 60411, 60411, 60411, 60411, 60411, 60411, 60411, 60386, 60386, 60386, 60386, 60386, 60386, 60355, 60355, 60355, 60355, 60355, 60355, 60355, 60330, 60330, 60330, 60330, 60330, 60330, 60330, 60298, 60298, 60298, 60298, 60298, 60298, 60273, 60273, 60273, 60273, 60273, 60273, 60273, 60242, 60242, 60242, 60242, 60242, 60242, 60242, 60217, 60217, 60217, 60217, 60217, 60217, 60185, 60185, 60185, 60185, 60185, 60185, 60185, 60160, 60160, 60160, 60160, 60160, 60160, 60129, 60129, 60129, 60129, 60129, 60129, 60129, 60104, 60104, 60104, 60104, 60104, 60104, 60104, 60073, 60073, 60073, 60073, 60073, 60073, 60048, 60048, 60048, 60048, 60048, 60048, 60048, 60017, 60017, 60017, 60017, 60017, 60017, 59992, 59992, 59992, 59992, 59992, 59992, 59992, 59960, 59960, 59960, 59960, 59960, 59960, 59960, 59935, 59935, 59935, 59935, 59935, 59935, 59910, 59910, 59910, 59910, 59910, 59910, 59910, 59879, 59879, 59879, 59879, 59879, 59879, 59854, 59854, 59854, 59854, 59854, 59854, 59854, 59823, 59823, 59823, 59823, 59823, 59823, 59798, 59798, 59798, 59798, 59798, 59798, 59798, 59767, 59767, 59767, 59767, 59767, 59767, 59742, 59742, 59742, 59742, 59742, 59742, 59742, 59711, 59711, 59711, 59711, 59711, 59711, 59686, 59686, 59686, 59686, 59686, 59686, 59686, 59655, 59655, 59655, 59655, 59655, 59655, 59630, 59630, 59630, 59630, 59630, 59630, 59630, 59599, 59599, 59599, 59599, 59599, 59599, 59574, 59574, 59574, 59574, 59574, 59574, 59574, 59543, 59543, 59543, 59543, 59543, 59543, 59518, 59518, 59518, 59518, 59518, 59518, 59518, 59487, 59487, 59487, 59487, 59487, 59487, 59462, 59462, 59462, 59462, 59462, 59462, 59431, 59431, 59431, 59431, 59431, 59431, 59431, 59406, 59406, 59406, 59406, 59406, 59406, 59375, 59375, 59375, 59375, 59375, 59375, 59375, 59350, 59350, 59350, 59350, 59350, 59350, 59319, 59319, 59319, 59319, 59319, 59319, 59295, 59295, 59295, 59295, 59295, 59295, 59295, 59264, 59264, 59264, 59264, 59264, 59264, 59239, 59239, 59239, 59239, 59239, 59239, 59239, 59208, 59208, 59208, 59208, 59208, 59208, 59183, 59183, 59183, 59183, 59183, 59183, 59152, 59152, 59152, 59152, 59152, 59152, 59152, 59127, 59127, 59127, 59127, 59127, 59127, 59096, 59096, 59096, 59096, 59096, 59096, 59072, 59072, 59072, 59072, 59072, 59072, 59072, 59041, 59041, 59041, 59041, 59041, 59041, 59016, 59016, 59016, 59016, 59016, 59016, 58985, 58985, 58985, 58985, 58985, 58985, 58985, 58960, 58960, 58960, 58960, 58960, 58960, 58929, 58929, 58929, 58929, 58929, 58929, 58905, 58905, 58905, 58905, 58905, 58905, 58905, 58874, 58874, 58874, 58874, 58874, 58874, 58849, 58849, 58849, 58849, 58849, 58849, 58818, 58818, 58818, 58818, 58818, 58818, 58794, 58794, 58794, 58794, 58794, 58794, 58794, 58763, 58763, 58763, 58763, 58763, 58763, 58738, 58738, 58738, 58738, 58738, 58738, 58707, 58707, 58707, 58707, 58707, 58707, 58683, 58683, 58683, 58683, 58683, 58683, 58683, 58658, 58658, 58658, 58658, 58658, 58658, 58627, 58627, 58627, 58627, 58627, 58627, 58603, 58603, 58603, 58603, 58603, 58603, 58572, 58572, 58572, 58572, 58572, 58572, 58547, 58547, 58547, 58547, 58547, 58547, 58547, 58516, 58516, 58516, 58516, 58516, 58516, 58492, 58492, 58492, 58492, 58492, 58492, 58461, 58461, 58461, 58461, 58461, 58461, 58436, 58436, 58436, 58436, 58436, 58436, 58406, 58406, 58406, 58406, 58406, 58406, 58406, 58381, 58381, 58381, 58381, 58381, 58381, 58350, 58350, 58350, 58350, 58350, 58350, 58326, 58326, 58326, 58326, 58326, 58326, 58295, 58295, 58295, 58295, 58295, 58295, 58271, 58271, 58271, 58271, 58271, 58271, 58240, 58240, 58240, 58240, 58240, 58240, 58215, 58215, 58215, 58215, 58215, 58215, 58215, 58185, 58185, 58185, 58185, 58185, 58185, 58160, 58160, 58160, 58160, 58160, 58160, 58130, 58130, 58130, 58130, 58130, 58130, 58105, 58105, 58105, 58105, 58105, 58105, 58075, 58075, 58075, 58075, 58075, 58075, 58050, 58050, 58050, 58050, 58050, 58050, 58019, 58019, 58019, 58019, 58019, 58019, 57995, 57995, 57995, 57995, 57995, 57995, 57964, 57964, 57964, 57964, 57964, 57964, 57940, 57940, 57940, 57940, 57940, 57940, 57940, 57909, 57909, 57909, 57909, 57909, 57909, 57885, 57885, 57885, 57885, 57885, 57885, 57854, 57854, 57854, 57854, 57854, 57854, 57830, 57830, 57830, 57830, 57830, 57830, 57799, 57799, 57799, 57799, 57799, 57799, 57775, 57775, 57775, 57775, 57775, 57775, 57744, 57744, 57744, 57744, 57744, 57744, 57720, 57720, 57720, 57720, 57720, 57720, 57689, 57689, 57689, 57689, 57689, 57689, 57665, 57665, 57665, 57665, 57665, 57665, 57635, 57635, 57635, 57635, 57635, 57635, 57610, 57610, 57610, 57610, 57610, 57610, 57580, 57580, 57580, 57580, 57580, 57580, 57555, 57555, 57555, 57555, 57555, 57555, 57525, 57525, 57525, 57525, 57525, 57525, 57501, 57501, 57501, 57501, 57501, 57501, 57470, 57470, 57470, 57470, 57470, 57470, 57446, 57446, 57446, 57446, 57446, 57446, 57421, 57421, 57421, 57421, 57421, 57421, 57391, 57391, 57391, 57391, 57391, 57391, 57367, 57367, 57367, 57367, 57367, 57367, 57336, 57336, 57336, 57336, 57336, 57312, 57312, 57312, 57312, 57312, 57312, 57282, 57282, 57282, 57282, 57282, 57282, 57257, 57257, 57257, 57257, 57257, 57257, 57227, 57227, 57227, 57227, 57227, 57227, 57203, 57203, 57203, 57203, 57203, 57203, 57172, 57172, 57172, 57172, 57172, 57172, 57148, 57148, 57148, 57148, 57148, 57148, 57118, 57118, 57118, 57118, 57118, 57118, 57093, 57093, 57093, 57093, 57093, 57093, 57063, 57063, 57063, 57063, 57063, 57063, 57039, 57039, 57039, 57039, 57039, 57009, 57009, 57009, 57009, 57009, 57009, 56984, 56984, 56984, 56984, 56984, 56984, 56954, 56954, 56954, 56954, 56954, 56954, 56930, 56930, 56930, 56930, 56930, 56930, 56900, 56900, 56900, 56900, 56900, 56900, 56875, 56875, 56875, 56875, 56875, 56875, 56845, 56845, 56845, 56845, 56845, 56821, 56821, 56821, 56821, 56821, 56821, 56791, 56791, 56791, 56791, 56791, 56791, 56767, 56767, 56767, 56767, 56767, 56767, 56736, 56736, 56736, 56736, 56736, 56736, 56712, 56712, 56712, 56712, 56712, 56712, 56682, 56682, 56682, 56682, 56682, 56658, 56658, 56658, 56658, 56658, 56658, 56628, 56628, 56628, 56628, 56628, 56628, 56603, 56603, 56603, 56603, 56603, 56603, 56573, 56573, 56573, 56573, 56573, 56573, 56549, 56549, 56549, 56549, 56549, 56519, 56519, 56519, 56519, 56519, 56519, 56495, 56495, 56495, 56495, 56495, 56495, 56465, 56465, 56465, 56465, 56465, 56465, 56441, 56441, 56441, 56441, 56441, 56410, 56410, 56410, 56410, 56410, 56410, 56386, 56386, 56386, 56386, 56386, 56386, 56356, 56356, 56356, 56356, 56356, 56356, 56332, 56332, 56332, 56332, 56332, 56302, 56302, 56302, 56302, 56302, 56302, 56278, 56278, 56278, 56278, 56278, 56278, 56254, 56254, 56254, 56254, 56254, 56254, 56224, 56224, 56224, 56224, 56224, 56200, 56200, 56200, 56200, 56200, 56200, 56170, 56170, 56170, 56170, 56170, 56170, 56146, 56146, 56146, 56146, 56146, 56116, 56116, 56116, 56116, 56116, 56116, 56092, 56092, 56092, 56092, 56092, 56092, 56062, 56062, 56062, 56062, 56062, 56062, 56038, 56038, 56038, 56038, 56038, 56008, 56008, 56008, 56008, 56008, 56008, 55984, 55984, 55984, 55984, 55984, 55984, 55954, 55954, 55954, 55954, 55954, 55930, 55930, 55930, 55930, 55930, 55930, 55900, 55900, 55900, 55900, 55900, 55900, 55876, 55876, 55876, 55876, 55876, 55846, 55846, 55846, 55846, 55846, 55846, 55822, 55822, 55822, 55822, 55822, 55822, 55792, 55792, 55792, 55792, 55792, 55768, 55768, 55768, 55768, 55768, 55768, 55738, 55738, 55738, 55738, 55738, 55714, 55714, 55714, 55714, 55714, 55714, 55684, 55684, 55684, 55684, 55684, 55684, 55660, 55660, 55660, 55660, 55660, 55630, 55630, 55630, 55630, 55630, 55630, 55606, 55606, 55606, 55606, 55606, 55606, 55576, 55576, 55576, 55576, 55576, 55552, 55552, 55552, 55552, 55552, 55552, 55523, 55523, 55523, 55523, 55523, 55499, 55499, 55499, 55499, 55499, 55499, 55469, 55469, 55469, 55469, 55469, 55469, 55445, 55445, 55445, 55445, 55445, 55415, 55415, 55415, 55415, 55415, 55415, 55391, 55391, 55391, 55391, 55391, 55361, 55361, 55361, 55361, 55361, 55361, 55338, 55338, 55338, 55338, 55338, 55308, 55308, 55308, 55308, 55308, 55308, 55284, 55284, 55284, 55284, 55284, 55284, 55254, 55254, 55254, 55254, 55254, 55230, 55230, 55230, 55230, 55230, 55230, 55200, 55200, 55200, 55200, 55200, 55177, 55177, 55177, 55177, 55177, 55177, 55147, 55147, 55147, 55147, 55147, 55123, 55123, 55123, 55123, 55123, 55123, 55093, 55093, 55093, 55093, 55093, 55069, 55069, 55069, 55069, 55069, 55069, 55046, 55046, 55046, 55046, 55046, 55016, 55016, 55016, 55016, 55016, 55016, 54992, 54992, 54992, 54992, 54992, 54962, 54962, 54962, 54962, 54962, 54962, 54939, 54939, 54939, 54939, 54939, 54909, 54909, 54909, 54909, 54909, 54909, 54885, 54885, 54885, 54885, 54885, 54855, 54855, 54855, 54855, 54855, 54855, 54832, 54832, 54832, 54832, 54832, 54802, 54802, 54802, 54802, 54802, 54802, 54778, 54778, 54778, 54778, 54778, 54749, 54749, 54749, 54749, 54749, 54749, 54725, 54725, 54725, 54725, 54725, 54695, 54695, 54695, 54695, 54695, 54695, 54671, 54671, 54671, 54671, 54671, 54642, 54642, 54642, 54642, 54642, 54642, 54618, 54618, 54618, 54618, 54618, 54588, 54588, 54588, 54588, 54588, 54565, 54565, 54565, 54565, 54565, 54565, 54535, 54535, 54535, 54535, 54535, 54511, 54511, 54511, 54511, 54511, 54511, 54482, 54482, 54482, 54482, 54482, 54458, 54458, 54458, 54458, 54458, 54458, 54429, 54429, 54429, 54429, 54429, 54405, 54405, 54405, 54405, 54405, 54375, 54375, 54375, 54375, 54375, 54375, 54352, 54352, 54352, 54352, 54352, 54322, 54322, 54322, 54322, 54322, 54322, 54299, 54299, 54299, 54299, 54299, 54269, 54269, 54269, 54269, 54269, 54245, 54245, 54245, 54245, 54245, 54245, 54216, 54216, 54216, 54216, 54216, 54192, 54192, 54192, 54192, 54192, 54192, 54163, 54163, 54163, 54163, 54163, 54139, 54139, 54139, 54139, 54139, 54110, 54110, 54110, 54110, 54110, 54110, 54086, 54086, 54086, 54086, 54086, 54056, 54056, 54056, 54056, 54056, 54033, 54033, 54033, 54033, 54033, 54033, 54003, 54003, 54003, 54003, 54003, 53980, 53980, 53980, 53980, 53980, 53950, 53950, 53950, 53950, 53950, 53950, 53927, 53927, 53927, 53927, 53927, 53897, 53897, 53897, 53897, 53897, 53897, 53874, 53874, 53874, 53874, 53874, 53850, 53850, 53850, 53850, 53850, 53821, 53821, 53821, 53821, 53821, 53821, 53797, 53797, 53797, 53797, 53797, 53768, 53768, 53768, 53768, 53768, 53744, 53744, 53744, 53744, 53744, 53715, 53715, 53715, 53715, 53715, 53715, 53691, 53691, 53691, 53691, 53691, 53662, 53662, 53662, 53662, 53662, 53638, 53638, 53638, 53638, 53638, 53638, 53609, 53609, 53609, 53609, 53609, 53586, 53586, 53586, 53586, 53586, 53556, 53556, 53556, 53556, 53556, 53556, 53533, 53533, 53533, 53533, 53533, 53503, 53503, 53503, 53503, 53503, 53480, 53480, 53480, 53480, 53480, 53451, 53451, 53451, 53451, 53451, 53451, 53427, 53427, 53427, 53427, 53427, 53398, 53398, 53398, 53398, 53398, 53374, 53374, 53374, 53374, 53374, 53345, 53345, 53345, 53345, 53345, 53345, 53322, 53322, 53322, 53322, 53322, 53292, 53292, 53292, 53292, 53292, 53269, 53269, 53269, 53269, 53269, 53240, 53240, 53240, 53240, 53240, 53240, 53216, 53216, 53216, 53216, 53216, 53187, 53187, 53187, 53187, 53187, 53163, 53163, 53163, 53163, 53163, 53134, 53134, 53134, 53134, 53134, 53134, 53111, 53111, 53111, 53111, 53111, 53081, 53081, 53081, 53081, 53081, 53058, 53058, 53058, 53058, 53058, 53029, 53029, 53029, 53029, 53029, 53029, 53005, 53005, 53005, 53005, 53005, 52976, 52976, 52976, 52976, 52976, 52953, 52953, 52953, 52953, 52953, 52924, 52924, 52924, 52924, 52924, 52900, 52900, 52900, 52900, 52900, 52900, 52871, 52871, 52871, 52871, 52871, 52848, 52848, 52848, 52848, 52848, 52819, 52819, 52819, 52819, 52819, 52795, 52795, 52795, 52795, 52795, 52766, 52766, 52766, 52766, 52766, 52743, 52743, 52743, 52743, 52743, 52743, 52713, 52713, 52713, 52713, 52713, 52690, 52690, 52690, 52690, 52690, 52667, 52667, 52667, 52667, 52667, 52638, 52638, 52638, 52638, 52638, 52614, 52614, 52614, 52614, 52614, 52585, 52585, 52585, 52585, 52585, 52585, 52562, 52562, 52562, 52562, 52562, 52533, 52533, 52533, 52533, 52533, 52510, 52510, 52510, 52510, 52510, 52480, 52480, 52480, 52480, 52480, 52457, 52457, 52457, 52457, 52457, 52428, 52428, 52428, 52428, 52428, 52405, 52405, 52405, 52405, 52405, 52405, 52376, 52376, 52376, 52376, 52376, 52352, 52352, 52352, 52352, 52352, 52323, 52323, 52323, 52323, 52323, 52300, 52300, 52300, 52300, 52300, 52271, 52271, 52271, 52271, 52271, 52248, 52248, 52248, 52248, 52248, 52219, 52219, 52219, 52219, 52219, 52195, 52195, 52195, 52195, 52195, 52195, 52166, 52166, 52166, 52166, 52166, 52143, 52143, 52143, 52143, 52143, 52114, 52114, 52114, 52114, 52114, 52091, 52091, 52091, 52091, 52091, 52062, 52062, 52062, 52062, 52062, 52039, 52039, 52039, 52039, 52039, 52010, 52010, 52010, 52010, 52010, 51987, 51987, 51987, 51987, 51987, 51958, 51958, 51958, 51958, 51958, 51934, 51934, 51934, 51934, 51934, 51905, 51905, 51905, 51905, 51905, 51882, 51882, 51882, 51882, 51882, 51853, 51853, 51853, 51853, 51853, 51853, 51830, 51830, 51830, 51830, 51830, 51801, 51801, 51801, 51801, 51801, 51778, 51778, 51778, 51778, 51778, 51749, 51749, 51749, 51749, 51749, 51726, 51726, 51726, 51726, 51726, 51697, 51697, 51697, 51697, 51697, 51674, 51674, 51674, 51674, 51674, 51645, 51645, 51645, 51645, 51645, 51622, 51622, 51622, 51622, 51622, 51593, 51593, 51593, 51593, 51593, 51570, 51570, 51570, 51570, 51570, 51547, 51547, 51547, 51547, 51547, 51518, 51518, 51518, 51518, 51518, 51495, 51495, 51495, 51495, 51495, 51466, 51466, 51466, 51466, 51466, 51443, 51443, 51443, 51443, 51443, 51414, 51414, 51414, 51414, 51414, 51391, 51391, 51391, 51391, 51391, 51362, 51362, 51362, 51362, 51362, 51339, 51339, 51339, 51339, 51339, 51310, 51310, 51310, 51310, 51310, 51287, 51287, 51287, 51287, 51287, 51258, 51258, 51258, 51258, 51258, 51235, 51235, 51235, 51235, 51235, 51206, 51206, 51206, 51206, 51206, 51183, 51183, 51183, 51183, 51183, 51154, 51154, 51154, 51154, 51154, 51131, 51131, 51131, 51131, 51131, 51102, 51102, 51102, 51102, 51102, 51079, 51079, 51079, 51079, 51079, 51050, 51050, 51050, 51050, 51050, 51027, 51027, 51027, 51027, 51027, 50999, 50999, 50999, 50999, 50999, 50976, 50976, 50976, 50976, 50976, 50947, 50947, 50947, 50947, 50947, 50924, 50924, 50924, 50924, 50924, 50895, 50895, 50895, 50895, 50872, 50872, 50872, 50872, 50872, 50843, 50843, 50843, 50843, 50843, 50820, 50820, 50820, 50820, 50820, 50792, 50792, 50792, 50792, 50792, 50769, 50769, 50769, 50769, 50769, 50740, 50740, 50740, 50740, 50740, 50717, 50717, 50717, 50717, 50717, 50688, 50688, 50688, 50688, 50688, 50665, 50665, 50665, 50665, 50665, 50636, 50636, 50636, 50636, 50636, 50613, 50613, 50613, 50613, 50613, 50585, 50585, 50585, 50585, 50585, 50562, 50562, 50562, 50562, 50533, 50533, 50533, 50533, 50533, 50510, 50510, 50510, 50510, 50510, 50482, 50482, 50482, 50482, 50482, 50459, 50459, 50459, 50459, 50459, 50430, 50430, 50430, 50430, 50430, 50407, 50407, 50407, 50407, 50407, 50384, 50384, 50384, 50384, 50384, 50355, 50355, 50355, 50355, 50355, 50332, 50332, 50332, 50332, 50304, 50304, 50304, 50304, 50304, 50281, 50281, 50281, 50281, 50281, 50252, 50252, 50252, 50252, 50252, 50229, 50229, 50229, 50229, 50229, 50201, 50201, 50201, 50201, 50201, 50178, 50178, 50178, 50178, 50178, 50149, 50149, 50149, 50149, 50149, 50126, 50126, 50126, 50126, 50098, 50098, 50098, 50098, 50098, 50075, 50075, 50075, 50075, 50075, 50046, 50046, 50046, 50046, 50046, 50023, 50023, 50023, 50023, 50023, 49995, 49995, 49995, 49995, 49995, 49972, 49972, 49972, 49972, 49943, 49943, 49943, 49943, 49943, 49921, 49921, 49921, 49921, 49921, 49892, 49892, 49892, 49892, 49892, 49869, 49869, 49869, 49869, 49869, 49841, 49841, 49841, 49841, 49841, 49818, 49818, 49818, 49818, 49789, 49789, 49789, 49789, 49789, 49766, 49766, 49766, 49766, 49766, 49738, 49738, 49738, 49738, 49738, 49715, 49715, 49715, 49715, 49715, 49687, 49687, 49687, 49687, 49687, 49664, 49664, 49664, 49664, 49635, 49635, 49635, 49635, 49635, 49612, 49612, 49612, 49612, 49612, 49584, 49584, 49584, 49584, 49584, 49561, 49561, 49561, 49561, 49561, 49533, 49533, 49533, 49533, 49510, 49510, 49510, 49510, 49510, 49481, 49481, 49481, 49481, 49481, 49459, 49459, 49459, 49459, 49459, 49430, 49430, 49430, 49430, 49407, 49407, 49407, 49407, 49407, 49379, 49379, 49379, 49379, 49379, 49356, 49356, 49356, 49356, 49356, 49328, 49328, 49328, 49328, 49328, 49305, 49305, 49305, 49305, 49276, 49276, 49276, 49276, 49276, 49254, 49254, 49254, 49254, 49254, 49231, 49231, 49231, 49231, 49231, 49203, 49203, 49203, 49203, 49180, 49180, 49180, 49180, 49180, 49151, 49151, 49151, 49151, 49151, 49129, 49129, 49129, 49129, 49129, 49100, 49100, 49100, 49100, 49078, 49078, 49078, 49078, 49078, 49049, 49049, 49049, 49049, 49049, 49026, 49026, 49026, 49026, 49026, 48998, 48998, 48998, 48998, 48975, 48975, 48975, 48975, 48975, 48947, 48947, 48947, 48947, 48947, 48924, 48924, 48924, 48924, 48924, 48896, 48896, 48896, 48896, 48873, 48873, 48873, 48873, 48873, 48845, 48845, 48845, 48845, 48845, 48822, 48822, 48822, 48822, 48794, 48794, 48794, 48794, 48794, 48771, 48771, 48771, 48771, 48771, 48743, 48743, 48743, 48743, 48743, 48720, 48720, 48720, 48720, 48692, 48692, 48692, 48692, 48692, 48669, 48669, 48669, 48669, 48669, 48641, 48641, 48641, 48641, 48618, 48618, 48618, 48618, 48618, 48590, 48590, 48590, 48590, 48590, 48567, 48567, 48567, 48567, 48539, 48539, 48539, 48539, 48539, 48516, 48516, 48516, 48516, 48516, 48488, 48488, 48488, 48488, 48488, 48465, 48465, 48465, 48465, 48437, 48437, 48437, 48437, 48437, 48414, 48414, 48414, 48414, 48414, 48386, 48386, 48386, 48386, 48363, 48363, 48363, 48363, 48363, 48335, 48335, 48335, 48335, 48335, 48312, 48312, 48312, 48312, 48284, 48284, 48284, 48284, 48284, 48262, 48262, 48262, 48262, 48262, 48233, 48233, 48233, 48233, 48211, 48211, 48211, 48211, 48211, 48182, 48182, 48182, 48182, 48182, 48160, 48160, 48160, 48160, 48132, 48132, 48132, 48132, 48132, 48109, 48109, 48109, 48109, 48109, 48086, 48086, 48086, 48086, 48058, 48058, 48058, 48058, 48058, 48036, 48036, 48036, 48036, 48007, 48007, 48007, 48007, 48007, 47985, 47985, 47985, 47985, 47985, 47957, 47957, 47957, 47957, 47934, 47934, 47934, 47934, 47934, 47906, 47906, 47906, 47906, 47906, 47883, 47883, 47883, 47883, 47855, 47855, 47855, 47855, 47855, 47833, 47833, 47833, 47833, 47833, 47804, 47804, 47804, 47804, 47782, 47782, 47782, 47782, 47782, 47754, 47754, 47754, 47754, 47731, 47731, 47731, 47731, 47731, 47703, 47703, 47703, 47703, 47703, 47680, 47680, 47680, 47680, 47652, 47652, 47652, 47652, 47652, 47630, 47630, 47630, 47630, 47602, 47602, 47602, 47602, 47602, 47579, 47579, 47579, 47579, 47579, 47551, 47551, 47551, 47551, 47528, 47528, 47528, 47528, 47528, 47500, 47500, 47500, 47500, 47478, 47478, 47478, 47478, 47478, 47450, 47450, 47450, 47450, 47450, 47427, 47427, 47427, 47427, 47399, 47399, 47399, 47399, 47399, 47377, 47377, 47377, 47377, 47348, 47348, 47348, 47348, 47348, 47326, 47326, 47326, 47326, 47298, 47298, 47298, 47298, 47298, 47275, 47275, 47275, 47275, 47275, 47247, 47247, 47247, 47247, 47225, 47225, 47225, 47225, 47225, 47197, 47197, 47197, 47197, 47174, 47174, 47174, 47174, 47174, 47146, 47146, 47146, 47146, 47124, 47124, 47124, 47124, 47124, 47096, 47096, 47096, 47096, 47096, 47073, 47073, 47073, 47073, 47045, 47045, 47045, 47045, 47045, 47023, 47023, 47023, 47023, 46995, 46995, 46995, 46995, 46995, 46972, 46972, 46972, 46972, 46950, 46950, 46950, 46950, 46950, 46922, 46922, 46922, 46922, 46899, 46899, 46899, 46899, 46899, 46871, 46871, 46871, 46871, 46849, 46849, 46849, 46849, 46849, 46821, 46821, 46821, 46821, 46821, 46798, 46798, 46798, 46798, 46770, 46770, 46770, 46770, 46770, 46748, 46748, 46748, 46748, 46720, 46720, 46720, 46720, 46720, 46698, 46698, 46698, 46698, 46670, 46670, 46670, 46670, 46670, 46647, 46647, 46647, 46647, 46619, 46619, 46619, 46619, 46619, 46597, 46597, 46597, 46597, 46569, 46569, 46569, 46569, 46569, 46546, 46546, 46546, 46546, 46518, 46518, 46518, 46518, 46518, 46496, 46496, 46496, 46496, 46468, 46468, 46468, 46468, 46468, 46446, 46446, 46446, 46446, 46418, 46418, 46418, 46418, 46418, 46395, 46395, 46395, 46395, 46367, 46367, 46367, 46367, 46367, 46345, 46345, 46345, 46345, 46317, 46317, 46317, 46317, 46317, 46295, 46295, 46295, 46295, 46267, 46267, 46267, 46267, 46267, 46244, 46244, 46244, 46244, 46216, 46216, 46216, 46216, 46216, 46194, 46194, 46194, 46194, 46166, 46166, 46166, 46166, 46166, 46144, 46144, 46144, 46144, 46116, 46116, 46116, 46116, 46116, 46094, 46094, 46094, 46094, 46066, 46066, 46066, 46066, 46043, 46043, 46043, 46043, 46043, 46015, 46015, 46015, 46015, 45993, 45993, 45993, 45993, 45993, 45965, 45965, 45965, 45965, 45943, 45943, 45943, 45943, 45943, 45915, 45915, 45915, 45915, 45893, 45893, 45893, 45893, 45893, 45870, 45870, 45870, 45870, 45842, 45842, 45842, 45842, 45842, 45820, 45820, 45820, 45820, 45792, 45792, 45792, 45792, 45770, 45770, 45770, 45770, 45770, 45742, 45742, 45742, 45742, 45720, 45720, 45720, 45720, 45720, 45692, 45692, 45692, 45692, 45670, 45670, 45670, 45670, 45670, 45642, 45642, 45642, 45642, 45619, 45619, 45619, 45619, 45592, 45592, 45592, 45592, 45592, 45569, 45569, 45569, 45569, 45541, 45541, 45541, 45541, 45541, 45519, 45519, 45519, 45519, 45491, 45491, 45491, 45491, 45491, 45469, 45469, 45469, 45469, 45441, 45441, 45441, 45441, 45419, 45419, 45419, 45419, 45419, 45391, 45391, 45391, 45391, 45369, 45369, 45369, 45369, 45369, 45341, 45341, 45341, 45341, 45319, 45319, 45319, 45319, 45291, 45291, 45291, 45291, 45291, 45269, 45269, 45269, 45269, 45241, 45241, 45241, 45241, 45241, 45219, 45219, 45219, 45219, 45191, 45191, 45191, 45191, 45169, 45169, 45169, 45169, 45169, 45141, 45141, 45141, 45141, 45119, 45119, 45119, 45119, 45119, 45091, 45091, 45091, 45091, 45069, 45069, 45069, 45069, 45041, 45041, 45041, 45041, 45041, 45019, 45019, 45019, 45019, 44991, 44991, 44991, 44991, 44991, 44969, 44969, 44969, 44969, 44941, 44941, 44941, 44941, 44919, 44919, 44919, 44919, 44919, 44891, 44891, 44891, 44891, 44869, 44869, 44869, 44869, 44841, 44841, 44841, 44841, 44841, 44819, 44819, 44819, 44819, 44791, 44791, 44791, 44791, 44791, 44769, 44769, 44769, 44769, 44747, 44747, 44747, 44747, 44719, 44719, 44719, 44719, 44719, 44697, 44697, 44697, 44697, 44669, 44669, 44669, 44669, 44647, 44647, 44647, 44647, 44647, 44619, 44619, 44619, 44619, 44597, 44597, 44597, 44597, 44569, 44569, 44569, 44569, 44569, 44547, 44547, 44547, 44547, 44519, 44519, 44519, 44519, 44497, 44497, 44497, 44497, 44497, 44469, 44469, 44469, 44469, 44447, 44447, 44447, 44447, 44419, 44419, 44419, 44419, 44419, 44397, 44397, 44397, 44397, 44370, 44370, 44370, 44370, 44347, 44347, 44347, 44347, 44347, 44320, 44320, 44320, 44320, 44298, 44298, 44298, 44298, 44270, 44270, 44270, 44270, 44270, 44248, 44248, 44248, 44248, 44220, 44220, 44220, 44220, 44198, 44198, 44198, 44198, 44198, 44170, 44170, 44170, 44170, 44148, 44148, 44148, 44148, 44120, 44120, 44120, 44120, 44120, 44098, 44098, 44098, 44098, 44071, 44071, 44071, 44071, 44049, 44049, 44049, 44049, 44049, 44021, 44021, 44021, 44021, 43999, 43999, 43999, 43999, 43971, 43971, 43971, 43971, 43971, 43949, 43949, 43949, 43949, 43921, 43921, 43921, 43921, 43899, 43899, 43899, 43899, 43872, 43872, 43872, 43872, 43872, 43849, 43849, 43849, 43849, 43822, 43822, 43822, 43822, 43800, 43800, 43800, 43800, 43800, 43772, 43772, 43772, 43772, 43750, 43750, 43750, 43750, 43722, 43722, 43722, 43722, 43700, 43700, 43700, 43700, 43700, 43673, 43673, 43673, 43673, 43651, 43651, 43651, 43651, 43628, 43628, 43628, 43628, 43628, 43601, 43601, 43601, 43601, 43579, 43579, 43579, 43579, 43551, 43551, 43551, 43551, 43529, 43529, 43529, 43529, 43529, 43501, 43501, 43501, 43501, 43479, 43479, 43479, 43479, 43452, 43452, 43452, 43452, 43430, 43430, 43430, 43430, 43430, 43402, 43402, 43402, 43402, 43380, 43380, 43380, 43380, 43352, 43352, 43352, 43352, 43352, 43330, 43330, 43330, 43330, 43303, 43303, 43303, 43303, 43281, 43281, 43281, 43281, 43253, 43253, 43253, 43253, 43253, 43231, 43231, 43231, 43231, 43204, 43204, 43204, 43204, 43182, 43182, 43182, 43182, 43154, 43154, 43154, 43154, 43154, 43132, 43132, 43132, 43132, 43104, 43104, 43104, 43104, 43082, 43082, 43082, 43082, 43055, 43055, 43055, 43055, 43033, 43033, 43033, 43033, 43033, 43005, 43005, 43005, 43005, 42983, 42983, 42983, 42983, 42956, 42956, 42956, 42956, 42934, 42934, 42934, 42934, 42934, 42906, 42906, 42906, 42906, 42884, 42884, 42884, 42884, 42856, 42856, 42856, 42856, 42834, 42834, 42834, 42834, 42834, 42807, 42807, 42807, 42807, 42785, 42785, 42785, 42785, 42757, 42757, 42757, 42757, 42735, 42735, 42735, 42735, 42708, 42708, 42708, 42708, 42708, 42686, 42686, 42686, 42686, 42658, 42658, 42658, 42658, 42636, 42636, 42636, 42636, 42609, 42609, 42609, 42609, 42587, 42587, 42587, 42587, 42587, 42559, 42559, 42559, 42559, 42537, 42537, 42537, 42537, 42515, 42515, 42515, 42515, 42488, 42488, 42488, 42488, 42466, 42466, 42466, 42466, 42466, 42438, 42438, 42438, 42438, 42416, 42416, 42416, 42416, 42389, 42389, 42389, 42389, 42367, 42367, 42367, 42367, 42339, 42339, 42339, 42339, 42339, 42317, 42317, 42317, 42317, 42290, 42290, 42290, 42290, 42268, 42268, 42268, 42268, 42240, 42240, 42240, 42240, 42218, 42218, 42218, 42218, 42218, 42191, 42191, 42191, 42191, 42169, 42169, 42169, 42169, 42141, 42141, 42141, 42141, 42119, 42119, 42119, 42119, 42092, 42092, 42092, 42092, 42070, 42070, 42070, 42070, 42070, 42042, 42042, 42042, 42042, 42020, 42020, 42020, 42020, 41993, 41993, 41993, 41993, 41971, 41971, 41971, 41971, 41944, 41944, 41944, 41944, 41922, 41922, 41922, 41922, 41922, 41894, 41894, 41894, 41894, 41872, 41872, 41872, 41872, 41845, 41845, 41845, 41845, 41823, 41823, 41823, 41823, 41795, 41795, 41795, 41795, 41773, 41773, 41773, 41773, 41773, 41746, 41746, 41746, 41746, 41724, 41724, 41724, 41724, 41697, 41697, 41697, 41697, 41675, 41675, 41675, 41675, 41647, 41647, 41647, 41647, 41625, 41625, 41625, 41625, 41598, 41598, 41598, 41598, 41598, 41576, 41576, 41576, 41576, 41548, 41548, 41548, 41548, 41527, 41527, 41527, 41527, 41499, 41499, 41499, 41499, 41477, 41477, 41477, 41477, 41455, 41455, 41455, 41455, 41428, 41428, 41428, 41428, 41428, 41406, 41406, 41406, 41406, 41378, 41378, 41378, 41378, 41357, 41357, 41357, 41357, 41329, 41329, 41329, 41329, 41307, 41307, 41307, 41307, 41280, 41280, 41280, 41280, 41258, 41258, 41258, 41258, 41231, 41231, 41231, 41231, 41209, 41209, 41209, 41209, 41209, 41181, 41181, 41181, 41181, 41159, 41159, 41159, 41159, 41132, 41132, 41132, 41132, 41110, 41110, 41110, 41110, 41083, 41083, 41083, 41083, 41061, 41061, 41061, 41061, 41033, 41033, 41033, 41033, 41011, 41011, 41011, 41011, 40984, 40984, 40984, 40984, 40984, 40962, 40962, 40962, 40962, 40935, 40935, 40935, 40935, 40913, 40913, 40913, 40913, 40885, 40885, 40885, 40885, 40864, 40864, 40864, 40864, 40836, 40836, 40836, 40836, 40814, 40814, 40814, 40814, 40787, 40787, 40787, 40787, 40765, 40765, 40765, 40765, 40738, 40738, 40738, 40738, 40738, 40716, 40716, 40716, 40716, 40688, 40688, 40688, 40688, 40667, 40667, 40667, 40667, 40639, 40639, 40639, 40639, 40617, 40617, 40617, 40617, 40590, 40590, 40590, 40590, 40568, 40568, 40568, 40568, 40541, 40541, 40541, 40541, 40519, 40519, 40519, 40519, 40491, 40491, 40491, 40491, 40470, 40470, 40470, 40470, 40442, 40442, 40442, 40442, 40420, 40420, 40420, 40420, 40420, 40393, 40393, 40393, 40393, 40371, 40371, 40371, 40371, 40349, 40349, 40349, 40349, 40322, 40322, 40322, 40322, 40300, 40300, 40300, 40300, 40273, 40273, 40273, 40273, 40251, 40251, 40251, 40251, 40224, 40224, 40224, 40224, 40202, 40202, 40202, 40202, 40174, 40174, 40174, 40174, 40152, 40152, 40152, 40152, 40125, 40125, 40125, 40125, 40103, 40103, 40103, 40103, 40076, 40076, 40076, 40076, 40054, 40054, 40054, 40054, 40027, 40027, 40027, 40027, 40005, 40005, 40005, 40005, 39978, 39978, 39978, 39978, 39956, 39956, 39956, 39956, 39956, 39928, 39928, 39928, 39928, 39907, 39907, 39907, 39907, 39879, 39879, 39879, 39879, 39857, 39857, 39857, 39857, 39830, 39830, 39830, 39830, 39808, 39808, 39808, 39808, 39781, 39781, 39781, 39781, 39759, 39759, 39759, 39759, 39732, 39732, 39732, 39732, 39710, 39710, 39710, 39710, 39683, 39683, 39683, 39683, 39661, 39661, 39661, 39661, 39634, 39634, 39634, 39634, 39612, 39612, 39612, 39612, 39584, 39584, 39584, 39584, 39563, 39563, 39563, 39563, 39535, 39535, 39535, 39535, 39513, 39513, 39513, 39513, 39486, 39486, 39486, 39486, 39464, 39464, 39464, 39464, 39437, 39437, 39437, 39437, 39415, 39415, 39415, 39415, 39388, 39388, 39388, 39388, 39366, 39366, 39366, 39366, 39339, 39339, 39339, 39339, 39317, 39317, 39317, 39317, 39290, 39290, 39290, 39290, 39268, 39268, 39268, 39268, 39246, 39246, 39246, 39246, 39219, 39219, 39219, 39219, 39197, 39197, 39197, 39197, 39170, 39170, 39170, 39170, 39148, 39148, 39148, 39148, 39121, 39121, 39121, 39121, 39099, 39099, 39099, 39099, 39071, 39071, 39071, 39071, 39050, 39050, 39050, 39050, 39022, 39022, 39022, 39022, 39001, 39001, 39001, 39001, 38973, 38973, 38973, 38973, 38951, 38951, 38951, 38951, 38924, 38924, 38924, 38924, 38902, 38902, 38902, 38902, 38875, 38875, 38875, 38875, 38853, 38853, 38853, 38853, 38826, 38826, 38826, 38826, 38804, 38804, 38804, 38804, 38777, 38777, 38777, 38777, 38755, 38755, 38755, 38755, 38728, 38728, 38728, 38728, 38706, 38706, 38706, 38706, 38679, 38679, 38679, 38679, 38657, 38657, 38657, 38657, 38630, 38630, 38630, 38630, 38608, 38608, 38608, 38608, 38581, 38581, 38581, 38581, 38559, 38559, 38559, 38559, 38532, 38532, 38532, 38532, 38510, 38510, 38510, 38483, 38483, 38483, 38483, 38461, 38461, 38461, 38461, 38434, 38434, 38434, 38434, 38412, 38412, 38412, 38412, 38384, 38384, 38384, 38384, 38363, 38363, 38363, 38363, 38335, 38335, 38335, 38335, 38314, 38314, 38314, 38314, 38286, 38286, 38286, 38286, 38265, 38265, 38265, 38265, 38237, 38237, 38237, 38237, 38216, 38216, 38216, 38216, 38188, 38188, 38188, 38188, 38167, 38167, 38167, 38167, 38145, 38145, 38145, 38145, 38118, 38118, 38118, 38118, 38096, 38096, 38096, 38096, 38068, 38068, 38068, 38068, 38047, 38047, 38047, 38019, 38019, 38019, 38019, 37998, 37998, 37998, 37998, 37970, 37970, 37970, 37970, 37949, 37949, 37949, 37949, 37921, 37921, 37921, 37921, 37900, 37900, 37900, 37900, 37872, 37872, 37872, 37872, 37851, 37851, 37851, 37851, 37823, 37823, 37823, 37823, 37802, 37802, 37802, 37802, 37774, 37774, 37774, 37774, 37753, 37753, 37753, 37753, 37725, 37725, 37725, 37725, 37704, 37704, 37704, 37676, 37676, 37676, 37676, 37655, 37655, 37655, 37655, 37627, 37627, 37627, 37627, 37606, 37606, 37606, 37606, 37578, 37578, 37578, 37578, 37557, 37557, 37557, 37557, 37529, 37529, 37529, 37529, 37508, 37508, 37508, 37508, 37480, 37480, 37480, 37480, 37459, 37459, 37459, 37459, 37431, 37431, 37431, 37410, 37410, 37410, 37410, 37382, 37382, 37382, 37382, 37361, 37361, 37361, 37361, 37333, 37333, 37333, 37333, 37312, 37312, 37312, 37312, 37284, 37284, 37284, 37284, 37263, 37263, 37263, 37263, 37235, 37235, 37235, 37235, 37214, 37214, 37214, 37214, 37186, 37186, 37186, 37165, 37165, 37165, 37165, 37137, 37137, 37137, 37137, 37116, 37116, 37116, 37116, 37088, 37088, 37088, 37088, 37067, 37067, 37067, 37067, 37045, 37045, 37045, 37045, 37018, 37018, 37018, 37018, 36996, 36996, 36996, 36969, 36969, 36969, 36969, 36947, 36947, 36947, 36947, 36920, 36920, 36920, 36920, 36898, 36898, 36898, 36898, 36871, 36871, 36871, 36871, 36849, 36849, 36849, 36849, 36822, 36822, 36822, 36822, 36800, 36800, 36800, 36800, 36773, 36773, 36773, 36751, 36751, 36751, 36751, 36724, 36724, 36724, 36724, 36702, 36702, 36702, 36702, 36675, 36675, 36675, 36675, 36653, 36653, 36653, 36653, 36626, 36626, 36626, 36626, 36604, 36604, 36604, 36577, 36577, 36577, 36577, 36555, 36555, 36555, 36555, 36528, 36528, 36528, 36528, 36506, 36506, 36506, 36506, 36479, 36479, 36479, 36479, 36457, 36457, 36457, 36457, 36430, 36430, 36430, 36408, 36408, 36408, 36408, 36381, 36381, 36381, 36381, 36359, 36359, 36359, 36359, 36332, 36332, 36332, 36332, 36310, 36310, 36310, 36310, 36283, 36283, 36283, 36283, 36261, 36261, 36261, 36234, 36234, 36234, 36234, 36212, 36212, 36212, 36212, 36185, 36185, 36185, 36185, 36163, 36163, 36163, 36163, 36136, 36136, 36136, 36136, 36114, 36114, 36114, 36087, 36087, 36087, 36087, 36065, 36065, 36065, 36065, 36038, 36038, 36038, 36038, 36016, 36016, 36016, 36016, 35995, 35995, 35995, 35995, 35967, 35967, 35967, 35946, 35946, 35946, 35946, 35918, 35918, 35918, 35918, 35897, 35897, 35897, 35897, 35869, 35869, 35869, 35869, 35848, 35848, 35848, 35848, 35820, 35820, 35820, 35799, 35799, 35799, 35799, 35771, 35771, 35771, 35771, 35750, 35750, 35750, 35750, 35722, 35722, 35722, 35722, 35701, 35701, 35701, 35701, 35674, 35674, 35674, 35652, 35652, 35652, 35652, 35625, 35625, 35625, 35625, 35603, 35603, 35603, 35603, 35576, 35576, 35576, 35576, 35554, 35554, 35554, 35527, 35527, 35527, 35527, 35505, 35505, 35505, 35505, 35478, 35478, 35478, 35478, 35456, 35456, 35456, 35456, 35429, 35429, 35429, 35407, 35407, 35407, 35407, 35380, 35380, 35380, 35380, 35358, 35358, 35358, 35358, 35331, 35331, 35331, 35331, 35309, 35309, 35309, 35309, 35282, 35282, 35282, 35260, 35260, 35260, 35260, 35233, 35233, 35233, 35233, 35211, 35211, 35211, 35211, 35184, 35184, 35184, 35184, 35162, 35162, 35162, 35135, 35135, 35135, 35135, 35113, 35113, 35113, 35113, 35086, 35086, 35086, 35086, 35064, 35064, 35064, 35037, 35037, 35037, 35037, 35015, 35015, 35015, 35015, 34988, 34988, 34988, 34988, 34966, 34966, 34966, 34966, 34939, 34939, 34939, 34917, 34917, 34917, 34917, 34895, 34895, 34895, 34895, 34868, 34868, 34868, 34868, 34846, 34846, 34846, 34846, 34819, 34819, 34819, 34797, 34797, 34797, 34797, 34770, 34770, 34770, 34770, 34748, 34748, 34748, 34748, 34721, 34721, 34721, 34699, 34699, 34699, 34699, 34672, 34672, 34672, 34672, 34650, 34650, 34650, 34650, 34623, 34623, 34623, 34623, 34601, 34601, 34601, 34574, 34574, 34574, 34574, 34552, 34552, 34552, 34552, 34525, 34525, 34525, 34525, 34503, 34503, 34503, 34476, 34476, 34476, 34476, 34454, 34454, 34454, 34454, 34427, 34427, 34427, 34427, 34405, 34405, 34405, 34378, 34378, 34378, 34378, 34356, 34356, 34356, 34356, 34329, 34329, 34329, 34329, 34307, 34307, 34307, 34280, 34280, 34280, 34280, 34258, 34258, 34258, 34258, 34231, 34231, 34231, 34231, 34209, 34209, 34209, 34182, 34182, 34182, 34182, 34160, 34160, 34160, 34160, 34133, 34133, 34133, 34133, 34111, 34111, 34111, 34084, 34084, 34084, 34084, 34062, 34062, 34062, 34062, 34035, 34035, 34035, 34035, 34013, 34013, 34013, 33986, 33986, 33986, 33986, 33964, 33964, 33964, 33964, 33937, 33937, 33937, 33937, 33915, 33915, 33915, 33888, 33888, 33888, 33888, 33866, 33866, 33866, 33866, 33839, 33839, 33839, 33839, 33817, 33817, 33817, 33795, 33795, 33795, 33795, 33768, 33768, 33768, 33768, 33746, 33746, 33746, 33746, 33719, 33719, 33719, 33697, 33697, 33697, 33697, 33670, 33670, 33670, 33670, 33648, 33648, 33648, 33648, 33621, 33621, 33621, 33599, 33599, 33599, 33599, 33572, 33572, 33572, 33572, 33550, 33550, 33550, 33523, 33523, 33523, 33523, 33501, 33501, 33501, 33501, 33474, 33474, 33474, 33474, 33452, 33452, 33452, 33425, 33425, 33425, 33425, 33403, 33403, 33403, 33403, 33376, 33376, 33376, 33354, 33354, 33354, 33354, 33327, 33327, 33327, 33327, 33305, 33305, 33305, 33305, 33278, 33278, 33278, 33256, 33256, 33256, 33256, 33229, 33229, 33229, 33229, 33207, 33207, 33207, 33179, 33179, 33179, 33179, 33158, 33158, 33158, 33158, 33130, 33130, 33130, 33130, 33109, 33109, 33109, 33081, 33081, 33081, 33081, 33059, 33059, 33059, 33059, 33032, 33032, 33032, 33010, 33010, 33010, 33010, 32983, 32983, 32983, 32983, 32961, 32961, 32961, 32961, 32934, 32934, 32934, 32912, 32912, 32912, 32912, 32885, 32885, 32885, 32885, 32863, 32863, 32863, 32836, 32836, 32836, 32836, 32814, 32814, 32814, 32814, 32787, 32787, 32787, 32765, 32765, 32765, 32765, 32738, 32738, 32738, 32738, 32716, 32716, 32716, 32716, 32694, 32694, 32694, 32667, 32667, 32667, 32667, 32645, 32645, 32645, 32645, 32618, 32618, 32618, 32596, 32596, 32596, 32596, 32568, 32568, 32568, 32568, 32547, 32547, 32547, 32519, 32519, 32519, 32519, 32498, 32498, 32498, 32498, 32470, 32470, 32470, 32448, 32448, 32448, 32448, 32421, 32421, 32421, 32421, 32399, 32399, 32399, 32372, 32372, 32372, 32372, 32350, 32350, 32350, 32350, 32323, 32323, 32323, 32301, 32301, 32301, 32301, 32274, 32274, 32274, 32274, 32252, 32252, 32252, 32225, 32225, 32225, 32225, 32203, 32203, 32203, 32203, 32175, 32175, 32175, 32154, 32154, 32154, 32154, 32126, 32126, 32126, 32126, 32104, 32104, 32104, 32077, 32077, 32077, 32077, 32055, 32055, 32055, 32055, 32028, 32028, 32028, 32006, 32006, 32006, 32006, 31979, 31979, 31979, 31979, 31957, 31957, 31957, 31930, 31930, 31930, 31930, 31908, 31908, 31908, 31908, 31880, 31880, 31880, 31858, 31858, 31858, 31858, 31831, 31831, 31831, 31831, 31809, 31809, 31809, 31782, 31782, 31782, 31782, 31760, 31760, 31760, 31760, 31733, 31733, 31733, 31711, 31711, 31711, 31711, 31684, 31684, 31684, 31684, 31662, 31662, 31662, 31640, 31640, 31640, 31640, 31612, 31612, 31612, 31612, 31591, 31591, 31591, 31563, 31563, 31563, 31563, 31541, 31541, 31541, 31541, 31514, 31514, 31514, 31492, 31492, 31492, 31492, 31465, 31465, 31465, 31465, 31443, 31443, 31443, 31416, 31416, 31416, 31416, 31394, 31394, 31394, 31366, 31366, 31366, 31366, 31344, 31344, 31344, 31344, 31317, 31317, 31317, 31295, 31295, 31295, 31295, 31268, 31268, 31268, 31268, 31246, 31246, 31246, 31219, 31219, 31219, 31219, 31197, 31197, 31197, 31197, 31169, 31169, 31169, 31147, 31147, 31147, 31147, 31120, 31120, 31120, 31098, 31098, 31098, 31098, 31071, 31071, 31071, 31071, 31049, 31049, 31049, 31021, 31021, 31021, 31021, 31000, 31000, 31000, 31000, 30972, 30972, 30972, 30950, 30950, 30950, 30950, 30923, 30923, 30923, 30901, 30901, 30901, 30901, 30874, 30874, 30874, 30874, 30852, 30852, 30852, 30824, 30824, 30824, 30824, 30802, 30802, 30802, 30802, 30775, 30775, 30775, 30753, 30753, 30753, 30753, 30726, 30726, 30726, 30704, 30704, 30704, 30704, 30676, 30676, 30676, 30676, 30654, 30654, 30654, 30627, 30627, 30627, 30627, 30605, 30605, 30605, 30605, 30578, 30578, 30578, 30556, 30556, 30556, 30556, 30534, 30534, 30534, 30506, 30506, 30506, 30506, 30484, 30484, 30484, 30484, 30457, 30457, 30457, 30435, 30435, 30435, 30435, 30408, 30408, 30408, 30386, 30386, 30386, 30386, 30358, 30358, 30358, 30358, 30336, 30336, 30336, 30309, 30309, 30309, 30309, 30287, 30287, 30287, 30260, 30260, 30260, 30260, 30238, 30238, 30238, 30238, 30210, 30210, 30210, 30188, 30188, 30188, 30188, 30161, 30161, 30161, 30139, 30139, 30139, 30139, 30111, 30111, 30111, 30111, 30089, 30089, 30089, 30062, 30062, 30062, 30062, 30040, 30040, 30040, 30012, 30012, 30012, 30012, 29991, 29991, 29991, 29991, 29963, 29963, 29963, 29941, 29941, 29941, 29941, 29914, 29914, 29914, 29892, 29892, 29892, 29892, 29864, 29864, 29864, 29842, 29842, 29842, 29842, 29815, 29815, 29815, 29815, 29793, 29793, 29793, 29765, 29765, 29765, 29765, 29743, 29743, 29743, 29716, 29716, 29716, 29716, 29694, 29694, 29694, 29694, 29666, 29666, 29666, 29644, 29644, 29644, 29644, 29617, 29617, 29617, 29595, 29595, 29595, 29595, 29567, 29567, 29567, 29545, 29545, 29545, 29545, 29518, 29518, 29518, 29518, 29496, 29496, 29496, 29468, 29468, 29468, 29468, 29446, 29446, 29446, 29424, 29424, 29424, 29424, 29397, 29397, 29397, 29375, 29375, 29375, 29375, 29347, 29347, 29347, 29347, 29325, 29325, 29325, 29298, 29298, 29298, 29298, 29276, 29276, 29276, 29248, 29248, 29248, 29248, 29226, 29226, 29226, 29199, 29199, 29199, 29199, 29177, 29177, 29177, 29177, 29149, 29149, 29149, 29127, 29127, 29127, 29127, 29100, 29100, 29100, 29078, 29078, 29078, 29078, 29050, 29050, 29050, 29028, 29028, 29028, 29028, 29000, 29000, 29000, 28978, 28978, 28978, 28978, 28951, 28951, 28951, 28951, 28929, 28929, 28929, 28901, 28901, 28901, 28901, 28879, 28879, 28879, 28852, 28852, 28852, 28852, 28830, 28830, 28830, 28802, 28802, 28802, 28802, 28780, 28780, 28780, 28752, 28752, 28752, 28752, 28730, 28730, 28730, 28730, 28703, 28703, 28703, 28681, 28681, 28681, 28681, 28653, 28653, 28653, 28631, 28631, 28631, 28631, 28603, 28603, 28603, 28581, 28581, 28581, 28581, 28554, 28554, 28554, 28532, 28532, 28532, 28532, 28504, 28504, 28504, 28482, 28482, 28482, 28482, 28454, 28454, 28454, 28454, 28432, 28432, 28432, 28405, 28405, 28405, 28405, 28383, 28383, 28383, 28355, 28355, 28355, 28355, 28333, 28333, 28333, 28311, 28311, 28311, 28311, 28283, 28283, 28283, 28261, 28261, 28261, 28261, 28233, 28233, 28233, 28211, 28211, 28211, 28211, 28184, 28184, 28184, 28162, 28162, 28162, 28162, 28134, 28134, 28134, 28112, 28112, 28112, 28112, 28084, 28084, 28084, 28084, 28062, 28062, 28062, 28034, 28034, 28034, 28034, 28012, 28012, 28012, 27985, 27985, 27985, 27985, 27963, 27963, 27963, 27935, 27935, 27935, 27935, 27913, 27913, 27913, 27885, 27885, 27885, 27885, 27863, 27863, 27863, 27835, 27835, 27835, 27835, 27813, 27813, 27813, 27785, 27785, 27785, 27785, 27763, 27763, 27763, 27736, 27736, 27736, 27736, 27713, 27713, 27713, 27686, 27686, 27686, 27686, 27664, 27664, 27664, 27636, 27636, 27636, 27636, 27614, 27614, 27614, 27586, 27586, 27586, 27586, 27564, 27564, 27564, 27536, 27536, 27536, 27536, 27514, 27514, 27514, 27486, 27486, 27486, 27486, 27464, 27464, 27464, 27436, 27436, 27436, 27436, 27414, 27414, 27414, 27387, 27387, 27387, 27387, 27364, 27364, 27364, 27337, 27337, 27337, 27337, 27314, 27314, 27314, 27287, 27287, 27287, 27287, 27264, 27264, 27264, 27237, 27237, 27237, 27237, 27215, 27215, 27215, 27192, 27192, 27192, 27192, 27165, 27165, 27165, 27142, 27142, 27142, 27142, 27115, 27115, 27115, 27092, 27092, 27092, 27092, 27065, 27065, 27065, 27042, 27042, 27042, 27042, 27015, 27015, 27015, 26992, 26992, 26992, 26992, 26965, 26965, 26965, 26942, 26942, 26942, 26942, 26915, 26915, 26915, 26892, 26892, 26892, 26892, 26865, 26865, 26865, 26842, 26842, 26842, 26842, 26815, 26815, 26815, 26792, 26792, 26792, 26792, 26765, 26765, 26765, 26742, 26742, 26742, 26742, 26715, 26715, 26715, 26692, 26692, 26692, 26692, 26664, 26664, 26664, 26642, 26642, 26642, 26642, 26614, 26614, 26614, 26592, 26592, 26592, 26592, 26564, 26564, 26564, 26542, 26542, 26542, 26542, 26514, 26514, 26514, 26492, 26492, 26492, 26492, 26464, 26464, 26464, 26442, 26442, 26442, 26442, 26414, 26414, 26414, 26392, 26392, 26392, 26392, 26364, 26364, 26364, 26342, 26342, 26342, 26342, 26314, 26314, 26314, 26291, 26291, 26291, 26264, 26264, 26264, 26264, 26241, 26241, 26241, 26213, 26213, 26213, 26213, 26191, 26191, 26191, 26163, 26163, 26163, 26163, 26141, 26141, 26141, 26119, 26119, 26119, 26119, 26091, 26091, 26091, 26068, 26068, 26068, 26068, 26040, 26040, 26040, 26018, 26018, 26018, 26018, 25990, 25990, 25990, 25968, 25968, 25968, 25968, 25940, 25940, 25940, 25918, 25918, 25918, 25890, 25890, 25890, 25890, 25867, 25867, 25867, 25839, 25839, 25839, 25839, 25817, 25817, 25817, 25789, 25789, 25789, 25789, 25767, 25767, 25767, 25739, 25739, 25739, 25739, 25717, 25717, 25717, 25689, 25689, 25689, 25689, 25666, 25666, 25666, 25638, 25638, 25638, 25638, 25616, 25616, 25616, 25588, 25588, 25588, 25566, 25566, 25566, 25566, 25538, 25538, 25538, 25515, 25515, 25515, 25515, 25487, 25487, 25487, 25465, 25465, 25465, 25465, 25437, 25437, 25437, 25414, 25414, 25414, 25414, 25386, 25386, 25386, 25364, 25364, 25364, 25336, 25336, 25336, 25336, 25314, 25314, 25314, 25286, 25286, 25286, 25286, 25263, 25263, 25263, 25235, 25235, 25235, 25235, 25213, 25213, 25213, 25185, 25185, 25185, 25185, 25162, 25162, 25162, 25134, 25134, 25134, 25112, 25112, 25112, 25112, 25084, 25084, 25084, 25061, 25061, 25061, 25061, 25033, 25033, 25033, 25011, 25011, 25011, 25011, 24989, 24989, 24989, 24960, 24960, 24960, 24960, 24938, 24938, 24938, 24910, 24910, 24910, 24887, 24887, 24887, 24887, 24859, 24859, 24859, 24837, 24837, 24837, 24837, 24809, 24809, 24809, 24786, 24786, 24786, 24786, 24758, 24758, 24758, 24736, 24736, 24736, 24708, 24708, 24708, 24708, 24685, 24685, 24685, 24657, 24657, 24657, 24657, 24635, 24635, 24635, 24607, 24607, 24607, 24607, 24584, 24584, 24584, 24556, 24556, 24556, 24533, 24533, 24533, 24533, 24505, 24505, 24505, 24483, 24483, 24483, 24483, 24455, 24455, 24455, 24432, 24432, 24432, 24432, 24404, 24404, 24404, 24381, 24381, 24381, 24353, 24353, 24353, 24353, 24331, 24331, 24331, 24303, 24303, 24303, 24303, 24280, 24280, 24280, 24252, 24252, 24252, 24229, 24229, 24229, 24229, 24201, 24201, 24201, 24179, 24179, 24179, 24179, 24150, 24150, 24150, 24128, 24128, 24128, 24128, 24100, 24100, 24100, 24077, 24077, 24077, 24049, 24049, 24049, 24049, 24026, 24026, 24026, 23998, 23998, 23998, 23998, 23976, 23976, 23976, 23947, 23947, 23947, 23925, 23925, 23925, 23925, 23897, 23897, 23897, 23874, 23874, 23874, 23874, 23851, 23851, 23851, 23823, 23823, 23823, 23801, 23801, 23801, 23801, 23772, 23772, 23772, 23750, 23750, 23750, 23750, 23721, 23721, 23721, 23699, 23699, 23699, 23671, 23671, 23671, 23671, 23648, 23648, 23648, 23620, 23620, 23620, 23620, 23597, 23597, 23597, 23569, 23569, 23569, 23546, 23546, 23546, 23546, 23518, 23518, 23518, 23495, 23495, 23495, 23495, 23467, 23467, 23467, 23444, 23444, 23444, 23416, 23416, 23416, 23416, 23393, 23393, 23393, 23365, 23365, 23365, 23365, 23342, 23342, 23342, 23314, 23314, 23314, 23291, 23291, 23291, 23291, 23263, 23263, 23263, 23240, 23240, 23240, 23240, 23212, 23212, 23212, 23189, 23189, 23189, 23161, 23161, 23161, 23161, 23138, 23138, 23138, 23110, 23110, 23110, 23110, 23087, 23087, 23087, 23059, 23059, 23059, 23036, 23036, 23036, 23036, 23008, 23008, 23008, 22985, 22985, 22985, 22957, 22957, 22957, 22957, 22934, 22934, 22934, 22905, 22905, 22905, 22905, 22883, 22883, 22883, 22854, 22854, 22854, 22832, 22832, 22832, 22832, 22803, 22803, 22803, 22780, 22780, 22780, 22752, 22752, 22752, 22752, 22729, 22729, 22729, 22706, 22706, 22706, 22706, 22678, 22678, 22678, 22655, 22655, 22655, 22627, 22627, 22627, 22627, 22604, 22604, 22604, 22576, 22576, 22576, 22576, 22553, 22553, 22553, 22524, 22524, 22524, 22502, 22502, 22502, 22502, 22473, 22473, 22473, 22450, 22450, 22450, 22422, 22422, 22422, 22422, 22399, 22399, 22399, 22370, 22370, 22370, 22348, 22348, 22348, 22348, 22319, 22319, 22319, 22296, 22296, 22296, 22296, 22268, 22268, 22268, 22245, 22245, 22245, 22216, 22216, 22216, 22216, 22194, 22194, 22194, 22165, 22165, 22165, 22142, 22142, 22142, 22142, 22114, 22114, 22114, 22091, 22091, 22091, 22062, 22062, 22062, 22062, 22039, 22039, 22039, 22011, 22011, 22011, 22011, 21988, 21988, 21988, 21959, 21959, 21959, 21937, 21937, 21937, 21937, 21908, 21908, 21908, 21885, 21885, 21885, 21856, 21856, 21856, 21856, 21834, 21834, 21834, 21805, 21805, 21805, 21782, 21782, 21782, 21782, 21753, 21753, 21753, 21731, 21731, 21731, 21731, 21702, 21702, 21702, 21679, 21679, 21679, 21650, 21650, 21650, 21650, 21627, 21627, 21627, 21604, 21604, 21604, 21576, 21576, 21576, 21576, 21553, 21553, 21553, 21524, 21524, 21524, 21501, 21501, 21501, 21501, 21473, 21473, 21473, 21450, 21450, 21450, 21421, 21421, 21421, 21421, 21398, 21398, 21398, 21369, 21369, 21369, 21346, 21346, 21346, 21346, 21318, 21318, 21318, 21295, 21295, 21295, 21266, 21266, 21266, 21266, 21243, 21243, 21243, 21214, 21214, 21214, 21191, 21191, 21191, 21191, 21162, 21162, 21162, 21139, 21139, 21139, 21111, 21111, 21111, 21111, 21088, 21088, 21088, 21059, 21059, 21059, 21036, 21036, 21036, 21036, 21007, 21007, 21007, 20984, 20984, 20984, 20984, 20955, 20955, 20955, 20932, 20932, 20932, 20904, 20904, 20904, 20904, 20880, 20880, 20880, 20852, 20852, 20852, 20829, 20829, 20829, 20829, 20800, 20800, 20800, 20777, 20777, 20777, 20748, 20748, 20748, 20748, 20725, 20725, 20725, 20696, 20696, 20696, 20673, 20673, 20673, 20644, 20644, 20644, 20644, 20621, 20621, 20621, 20592, 20592, 20592, 20569, 20569, 20569, 20569, 20540, 20540, 20540, 20517, 20517, 20517, 20488, 20488, 20488, 20488, 20465, 20465, 20465, 20442, 20442, 20442, 20413, 20413, 20413, 20413, 20390, 20390, 20390, 20361, 20361, 20361, 20338, 20338, 20338, 20338, 20309, 20309, 20309, 20286, 20286, 20286, 20257, 20257, 20257, 20257, 20234, 20234, 20234, 20205, 20205, 20205, 20182, 20182, 20182, 20182, 20153, 20153, 20153, 20129, 20129, 20129, 20100, 20100, 20100, 20100, 20077, 20077, 20077, 20048, 20048, 20048, 20025, 20025, 20025, 20025, 19996, 19996, 19996, 19973, 19973, 19973, 19944, 19944, 19944, 19921, 19921, 19921, 19921, 19892, 19892, 19892, 19868, 19868, 19868, 19839, 19839, 19839, 19839, 19816, 19816, 19816, 19787, 19787, 19787, 19764, 19764, 19764, 19764, 19735, 19735, 19735, 19712, 19712, 19712, 19682, 19682, 19682, 19682, 19659, 19659, 19659, 19630, 19630, 19630, 19607, 19607, 19607, 19607, 19578, 19578, 19578, 19555, 19555, 19555, 19525, 19525, 19525, 19502, 19502, 19502, 19502, 19473, 19473, 19473, 19450, 19450, 19450, 19421, 19421, 19421, 19421, 19397, 19397, 19397, 19368, 19368, 19368, 19345, 19345, 19345, 19345, 19316, 19316, 19316, 19292, 19292, 19292, 19269, 19269, 19269, 19240, 19240, 19240, 19240, 19217, 19217, 19217, 19187, 19187, 19187, 19164, 19164, 19164, 19164, 19135, 19135, 19135, 19111, 19111, 19111, 19082, 19082, 19082, 19082, 19059, 19059, 19059, 19030, 19030, 19030, 19006, 19006, 19006, 18977, 18977, 18977, 18977, 18954, 18954, 18954, 18924, 18924, 18924, 18901, 18901, 18901, 18901, 18872, 18872, 18872, 18848, 18848, 18848, 18819, 18819, 18819, 18796, 18796, 18796, 18796, 18766, 18766, 18766, 18743, 18743, 18743, 18714, 18714, 18714, 18714, 18690, 18690, 18690, 18661, 18661, 18661, 18637, 18637, 18637, 18608, 18608, 18608, 18608, 18585, 18585, 18585, 18555, 18555, 18555, 18532, 18532, 18532, 18532, 18502, 18502, 18502, 18479, 18479, 18479, 18450, 18450, 18450, 18426, 18426, 18426, 18426, 18397, 18397, 18397, 18373, 18373, 18373, 18344, 18344, 18344, 18344, 18320, 18320, 18320, 18291, 18291, 18291, 18267, 18267, 18267, 18238, 18238, 18238, 18238, 18215, 18215, 18215, 18185, 18185, 18185, 18162, 18162, 18162, 18162, 18132, 18132, 18132, 18109, 18109, 18109, 18085, 18085, 18085, 18056, 18056, 18056, 18056, 18032, 18032, 18032, 18002, 18002, 18002, 17979, 17979, 17979, 17949, 17949, 17949, 17949, 17926, 17926, 17926, 17896, 17896, 17896, 17873, 17873, 17873, 17873, 17843, 17843, 17843, 17820, 17820, 17820, 17790, 17790, 17790, 17766, 17766, 17766, 17766, 17737, 17737, 17737, 17713, 17713, 17713, 17684, 17684, 17684, 17660, 17660, 17660, 17660, 17631, 17631, 17631, 17607, 17607, 17607, 17577, 17577, 17577, 17554, 17554, 17554, 17554, 17524, 17524, 17524, 17500, 17500, 17500, 17471, 17471, 17471, 17471, 17447, 17447, 17447, 17417, 17417, 17417, 17394, 17394, 17394, 17364, 17364, 17364, 17364, 17340, 17340, 17340, 17311, 17311, 17311, 17287, 17287, 17287, 17257, 17257, 17257, 17257, 17234, 17234, 17234, 17204, 17204, 17204, 17180, 17180, 17180, 17151, 17151, 17151, 17151, 17127, 17127, 17127, 17097, 17097, 17097, 17073, 17073, 17073, 17044, 17044, 17044, 17044, 17020, 17020, 17020, 16990, 16990, 16990, 16966, 16966, 16966, 16937, 16937, 16937, 16937, 16913, 16913, 16913, 16889, 16889, 16889, 16859, 16859, 16859, 16835, 16835, 16835, 16835, 16806, 16806, 16806, 16782, 16782, 16782, 16752, 16752, 16752, 16728, 16728, 16728, 16728, 16698, 16698, 16698, 16674, 16674, 16674, 16645, 16645, 16645, 16621, 16621, 16621, 16621, 16591, 16591, 16591, 16567, 16567, 16567, 16537, 16537, 16537, 16513, 16513, 16513, 16513, 16483, 16483, 16483, 16459, 16459, 16459, 16430, 16430, 16430, 16406, 16406, 16406, 16406, 16376, 16376, 16376, 16352, 16352, 16352, 16322, 16322, 16322, 16298, 16298, 16298, 16298, 16268, 16268, 16268, 16244, 16244, 16244, 16214, 16214, 16214, 16190, 16190, 16190, 16190, 16160, 16160, 16160, 16136, 16136, 16136, 16106, 16106, 16106, 16082, 16082, 16082, 16082, 16052, 16052, 16052, 16028, 16028, 16028, 15998, 15998, 15998, 15974, 15974, 15974, 15944, 15944, 15944, 15944, 15920, 15920, 15920, 15890, 15890, 15890, 15866, 15866, 15866, 15836, 15836, 15836, 15836, 15812, 15812, 15812, 15782, 15782, 15782, 15758, 15758, 15758, 15734, 15734, 15734, 15734, 15704, 15704, 15704, 15680, 15680, 15680, 15650, 15650, 15650, 15626, 15626, 15626, 15596, 15596, 15596, 15596, 15571, 15571, 15571, 15541, 15541, 15541, 15517, 15517, 15517, 15487, 15487, 15487, 15487, 15463, 15463, 15463, 15433, 15433, 15433, 15409, 15409, 15409, 15378, 15378, 15378, 15378, 15354, 15354, 15354, 15324, 15324, 15324, 15300, 15300, 15300, 15270, 15270, 15270, 15246, 15246, 15246, 15246, 15215, 15215, 15215, 15191, 15191, 15191, 15161, 15161, 15161, 15137, 15137, 15137, 15137, 15106, 15106, 15106, 15082, 15082, 15082, 15052, 15052, 15052, 15028, 15028, 15028, 14997, 14997, 14997, 14997, 14973, 14973, 14973, 14943, 14943, 14943, 14919, 14919, 14919, 14888, 14888, 14888, 14864, 14864, 14864, 14864, 14834, 14834, 14834, 14809, 14809, 14809, 14779, 14779, 14779, 14755, 14755, 14755, 14755, 14724, 14724, 14724, 14700, 14700, 14700, 14670, 14670, 14670, 14645, 14645, 14645, 14615, 14615, 14615, 14615, 14591, 14591, 14591, 14560, 14560, 14560, 14536, 14536, 14536, 14512, 14512, 14512, 14481, 14481, 14481, 14481, 14457, 14457, 14457, 14426, 14426, 14426, 14402, 14402, 14402, 14371, 14371, 14371, 14371, 14347, 14347, 14347, 14317, 14317, 14317, 14292, 14292, 14292, 14262, 14262, 14262, 14237, 14237, 14237, 14237, 14207, 14207, 14207, 14182, 14182, 14182, 14152, 14152, 14152, 14127, 14127, 14127, 14097, 14097, 14097, 14097, 14072, 14072, 14072, 14042, 14042, 14042, 14017, 14017, 14017, 13987, 13987, 13987, 13962, 13962, 13962, 13962, 13932, 13932, 13932, 13907, 13907, 13907, 13876, 13876, 13876, 13852, 13852, 13852, 13821, 13821, 13821, 13821, 13797, 13797, 13797, 13766, 13766, 13766, 13742, 13742, 13742, 13711, 13711, 13711, 13686, 13686, 13686, 13686, 13656, 13656, 13656, 13631, 13631, 13631, 13600, 13600, 13600, 13576, 13576, 13576, 13545, 13545, 13545, 13545, 13521, 13521, 13521, 13490, 13490, 13490, 13465, 13465, 13465, 13434, 13434, 13434, 13410, 13410, 13410, 13379, 13379, 13379, 13379, 13354, 13354, 13354, 13324, 13324, 13324, 13299, 13299, 13299, 13274, 13274, 13274, 13243, 13243, 13243, 13243, 13219, 13219, 13219, 13188, 13188, 13188, 13163, 13163, 13163, 13132, 13132, 13132, 13108, 13108, 13108, 13108, 13077, 13077, 13077, 13052, 13052, 13052, 13021, 13021, 13021, 12996, 12996, 12996, 12966, 12966, 12966, 12941, 12941, 12941, 12941, 12910, 12910, 12910, 12885, 12885, 12885, 12854, 12854, 12854, 12829, 12829, 12829, 12798, 12798, 12798, 12798, 12774, 12774, 12774, 12743, 12743, 12743, 12718, 12718, 12718, 12687, 12687, 12687, 12662, 12662, 12662, 12631, 12631, 12631, 12631, 12606, 12606, 12606, 12575, 12575, 12575, 12550, 12550, 12550, 12519, 12519, 12519, 12494, 12494, 12494, 12494, 12463, 12463, 12463, 12438, 12438, 12438, 12407, 12407, 12407, 12382, 12382, 12382, 12351, 12351, 12351, 12326, 12326, 12326, 12326, 12295, 12295, 12295, 12270, 12270, 12270, 12239, 12239, 12239, 12214, 12214, 12214, 12183, 12183, 12183, 12158, 12158, 12158, 12158, 12127, 12127, 12127, 12102, 12102, 12102, 12071, 12071, 12071, 12046, 12046, 12046, 12021, 12021, 12021, 12021, 11990, 11990, 11990, 11965, 11965, 11965, 11933, 11933, 11933, 11908, 11908, 11908, 11877, 11877, 11877, 11852, 11852, 11852, 11852, 11821, 11821, 11821, 11796, 11796, 11796, 11764, 11764, 11764, 11739, 11739, 11739, 11708, 11708, 11708, 11683, 11683, 11683, 11683, 11652, 11652, 11652, 11627, 11627, 11627, 11595, 11595, 11595, 11570, 11570, 11570, 11539, 11539, 11539, 11514, 11514, 11514, 11514, 11482, 11482, 11482, 11457, 11457, 11457, 11426, 11426, 11426, 11400, 11400, 11400, 11369, 11369, 11369, 11344, 11344, 11344, 11312, 11312, 11312, 11312, 11287, 11287, 11287, 11256, 11256, 11256, 11231, 11231, 11231, 11199, 11199, 11199, 11174, 11174, 11174, 11142, 11142, 11142, 11142, 11117, 11117, 11117, 11085, 11085, 11085, 11060, 11060, 11060, 11029, 11029, 11029, 11003, 11003, 11003, 10972, 10972, 10972, 10972, 10947, 10947, 10947, 10915, 10915, 10915, 10890, 10890, 10890, 10858, 10858, 10858, 10833, 10833, 10833, 10807, 10807, 10807, 10776, 10776, 10776, 10776, 10750, 10750, 10750, 10719, 10719, 10719, 10693, 10693, 10693, 10662, 10662, 10662, 10636, 10636, 10636, 10605, 10605, 10605, 10579, 10579, 10579, 10579, 10548, 10548, 10548, 10522, 10522, 10522, 10490, 10490, 10490, 10465, 10465, 10465, 10433, 10433, 10433, 10408, 10408, 10408, 10408, 10376, 10376, 10376, 10351, 10351, 10351, 10319, 10319, 10319, 10293, 10293, 10293, 10261, 10261, 10261, 10236, 10236, 10236, 10204, 10204, 10204, 10204, 10179, 10179, 10179, 10147, 10147, 10147, 10121, 10121, 10121, 10089, 10089, 10089, 10064, 10064, 10064, 10032, 10032, 10032, 10006, 10006, 10006, 10006, 9974, 9974, 9974, 9949, 9949, 9949, 9917, 9917, 9917, 9891, 9891, 9891, 9859, 9859, 9859, 9834, 9834, 9834, 9802, 9802, 9802, 9802, 9776, 9776, 9776, 9744, 9744, 9744, 9718, 9718, 9718, 9686, 9686, 9686, 9661, 9661, 9661, 9629, 9629, 9629, 9603, 9603, 9603, 9571, 9571, 9571, 9571, 9545, 9545, 9545, 9520, 9520, 9520, 9487, 9487, 9487, 9462, 9462, 9462, 9430, 9430, 9430, 9404, 9404, 9404, 9372, 9372, 9372, 9372, 9346, 9346, 9346, 9314, 9314, 9314, 9288, 9288, 9288, 9256, 9256, 9256, 9230, 9230, 9230, 9198, 9198, 9198, 9172, 9172, 9172, 9140, 9140, 9140, 9140, 9114, 9114, 9114, 9082, 9082, 9082, 9056, 9056, 9056, 9024, 9024, 9024, 8998, 8998, 8998, 8965, 8965, 8965, 8940, 8940, 8940, 8907, 8907, 8907, 8907, 8881, 8881, 8881, 8849, 8849, 8849, 8823, 8823, 8823, 8791, 8791, 8791, 8765, 8765, 8765, 8732, 8732, 8732, 8706, 8706, 8706, 8674, 8674, 8674, 8674, 8648, 8648, 8648, 8616, 8616, 8616, 8590, 8590, 8590, 8557, 8557, 8557, 8531, 8531, 8531, 8499, 8499, 8499, 8473, 8473, 8473, 8440, 8440, 8440, 8440, 8414, 8414, 8414, 8382, 8382, 8382, 8356, 8356, 8356, 8323, 8323, 8323, 8297, 8297, 8297, 8264, 8264, 8264, 8238, 8238, 8238, 8212, 8212, 8212, 8212, 8180, 8180, 8180, 8153, 8153, 8153, 8121, 8121, 8121, 8095, 8095, 8095, 8062, 8062, 8062, 8036, 8036, 8036, 8003, 8003, 8003, 7977, 7977, 7977, 7944, 7944, 7944, 7944, 7918, 7918, 7918, 7885, 7885, 7885, 7859, 7859, 7859, 7827, 7827, 7827, 7800, 7800, 7800, 7768, 7768, 7768, 7741, 7741, 7741, 7708, 7708, 7708, 7682, 7682, 7682, 7682, 7649, 7649, 7649, 7623, 7623, 7623, 7590, 7590, 7590, 7564, 7564, 7564, 7531, 7531, 7531, 7505, 7505, 7505, 7472, 7472, 7472, 7446, 7446, 7446, 7413, 7413, 7413, 7413, 7386, 7386, 7386, 7353, 7353, 7353, 7327, 7327, 7327, 7294, 7294, 7294, 7268, 7268, 7268, 7235, 7235, 7235, 7208, 7208, 7208, 7175, 7175, 7175, 7149, 7149, 7149, 7149, 7116, 7116, 7116, 7089, 7089, 7089, 7056, 7056, 7056, 7030, 7030, 7030, 6997, 6997, 6997, 6970, 6970, 6970, 6937, 6937, 6937, 6911, 6911, 6911, 6884, 6884, 6884, 6851, 6851, 6851, 6851, 6825, 6825, 6825, 6791, 6791, 6791, 6765, 6765, 6765, 6732, 6732, 6732, 6705, 6705, 6705, 6672, 6672, 6672, 6645, 6645, 6645, 6612, 6612, 6612, 6585, 6585, 6585, 6552, 6552, 6552, 6552, 6525, 6525, 6525, 6492, 6492, 6492, 6466, 6466, 6466, 6432, 6432, 6432, 6406, 6406, 6406, 6372, 6372, 6372, 6346, 6346, 6346, 6312, 6312, 6312, 6285, 6285, 6285, 6252, 6252, 6252, 6252, 6225, 6225, 6225, 6192, 6192, 6192, 6165, 6165, 6165, 6132, 6132, 6132, 6105, 6105, 6105, 6072, 6072, 6072, 6045, 6045, 6045, 6011, 6011, 6011, 5984, 5984, 5984, 5951, 5951, 5951, 5924, 5924, 5924, 5924, 5891, 5891, 5891, 5864, 5864, 5864, 5830, 5830, 5830, 5803, 5803, 5803, 5770, 5770, 5770, 5743, 5743, 5743, 5709, 5709, 5709, 5682, 5682, 5682, 5649, 5649, 5649, 5622, 5622, 5622, 5588, 5588, 5588, 5561, 5561, 5561, 5561, 5534, 5534, 5534, 5500, 5500, 5500, 5473, 5473, 5473, 5440, 5440, 5440, 5413, 5413, 5413, 5379, 5379, 5379, 5352, 5352, 5352, 5318, 5318, 5318, 5291, 5291, 5291, 5257, 5257, 5257, 5230, 5230, 5230, 5196, 5196, 5196, 5196, 5169, 5169, 5169, 5135, 5135, 5135, 5108, 5108, 5108, 5074, 5074, 5074, 5047, 5047, 5047, 5013, 5013, 5013, 4986, 4986, 4986, 4952, 4952, 4952, 4925, 4925, 4925, 4891, 4891, 4891, 4864, 4864, 4864, 4830, 4830, 4830, 4830, 4803, 4803, 4803, 4769, 4769, 4769, 4741, 4741, 4741, 4707, 4707, 4707, 4680, 4680, 4680, 4646, 4646, 4646, 4619, 4619, 4619, 4585, 4585, 4585, 4557, 4557, 4557, 4523, 4523, 4523, 4496, 4496, 4496, 4462, 4462, 4462, 4434, 4434, 4434, 4434, 4400, 4400, 4400, 4373, 4373, 4373, 4339, 4339, 4339, 4311, 4311, 4311, 4277, 4277, 4277, 4250, 4250, 4250, 4222, 4222, 4222, 4188, 4188, 4188, 4161, 4161, 4161, 4126, 4126, 4126, 4099, 4099, 4099, 4064, 4064, 4064, 4037, 4037, 4037, 4003, 4003, 4003, 4003, 3975, 3975, 3975, 3941, 3941, 3941, 3913, 3913, 3913, 3879, 3879, 3879, 3851, 3851, 3851, 3817, 3817, 3817, 3789, 3789, 3789, 3755, 3755, 3755, 3727, 3727, 3727, 3693, 3693, 3693, 3665, 3665, 3665, 3631, 3631, 3631, 3603, 3603, 3603, 3568, 3568, 3568, 3541, 3541, 3541, 3541, 3506, 3506, 3506, 3478, 3478, 3478, 3444, 3444, 3444, 3416, 3416, 3416, 3381, 3381, 3381, 3354, 3354, 3354, 3319, 3319, 3319, 3291, 3291, 3291, 3257, 3257, 3257, 3229, 3229, 3229, 3194, 3194, 3194, 3166, 3166, 3166, 3132, 3132, 3132, 3104, 3104, 3104, 3069, 3069, 3069, 3041, 3041, 3041, 3041, 3006, 3006, 3006, 2978, 2978, 2978, 2944, 2944, 2944, 2916, 2916, 2916, 2881, 2881, 2881, 2853, 2853, 2853, 2825, 2825, 2825, 2790, 2790, 2790, 2762, 2762, 2762, 2727, 2727, 2727, 2699, 2699, 2699, 2664, 2664, 2664, 2636, 2636, 2636, 2601, 2601, 2601, 2573, 2573, 2573, 2538, 2538, 2538, 2510, 2510, 2510, 2475, 2475, 2475, 2475, 2447, 2447, 2447, 2412, 2412, 2412, 2384, 2384, 2384, 2349, 2349, 2349, 2321, 2321, 2321, 2285, 2285, 2285, 2257, 2257, 2257, 2222, 2222, 2222, 2194, 2194, 2194, 2159, 2159, 2159, 2131, 2131, 2131, 2095, 2095, 2095, 2067, 2067, 2067, 2032, 2032, 2032, 2004, 2004, 2004, 1968, 1968, 1968, 1940, 1940, 1940, 1905, 1905, 1905, 1876, 1876, 1876, 1841, 1841, 1841, 1841, 1813, 1813, 1813, 1777, 1777, 1777, 1749, 1749, 1749, 1714, 1714, 1714, 1685, 1685, 1685, 1650, 1650, 1650, 1621, 1621, 1621, 1586, 1586, 1586, 1558, 1558, 1558, 1522, 1522, 1522, 1494, 1494, 1494, 1458, 1458, 1458, 1430, 1430, 1430, 1401, 1401, 1401, 1366, 1366, 1366, 1337, 1337, 1337, 1301, 1301, 1301, 1273, 1273, 1273, 1237, 1237, 1237, 1209, 1209, 1209, 1173, 1173, 1173, 1144, 1144, 1144, 1144, 1109, 1109, 1109, 1080, 1080, 1080, 1044, 1044, 1044, 1016, 1016, 1016, 980, 980, 980, 951, 951, 951, 916, 916, 916, 887, 887, 887, 851, 851, 851, 822, 822, 822, 787, 787, 787, 758, 758, 758, 722, 722, 722, 693, 693, 693, 657, 657, 657, 628, 628, 628, 592, 592, 592, 564, 564, 564, 528, 528, 528, 499, 499, 499, 463, 463, 463, 434, 434, 434, 398, 398, 398, 369, 369, 369, 333, 333, 333, 304, 304, 304, 268, 268, 268, 268, 239, 239, 239, 203, 203, 203, 174, 174, 174, 138, 138, 138, 109, 109, 109, 73, 73, 73, 44, 44, 44, 7, 7, 7, 71978, 71978, 71978, 71949, 71949, 71949, 71913, 71913, 71913, 71884, 71884, 71884, 71848, 71848, 71848, 71819, 71819, 71819, 71783, 71783, 71783, 71754, 71754, 71754, 71718, 71718, 71718, 71689, 71689, 71689, 71653, 71653, 71653, 71624, 71624, 71624, 71588, 71588, 71588, 71559, 71559, 71559, 71523, 71523, 71523, 71494, 71494, 71494, 71458, 71458, 71458, 71429, 71429, 71429, 71393, 71393, 71393, 71364, 71364, 71364, 71328, 71328, 71328, 71300, 71300, 71300, 71264, 71264, 71264, 71235, 71235, 71235, 71199, 71199, 71199, 71170, 71170, 71170, 71135, 71135, 71135, 71106, 71106, 71106, 71106, 71070, 71070, 71070, 71041, 71041, 71041, 71006, 71006, 71006, 70977, 70977, 70977, 70941, 70941, 70941, 70913, 70913, 70913, 70877, 70877, 70877, 70848, 70848, 70848, 70813, 70813, 70813, 70784, 70784, 70784, 70748, 70748, 70748, 70720, 70720, 70720, 70684, 70684, 70684, 70656, 70656, 70656, 70620, 70620, 70620, 70592, 70592, 70592, 70563, 70563, 70563, 70528, 70528, 70528, 70499, 70499, 70499, 70464, 70464, 70464, 70435, 70435, 70435, 70400, 70400, 70400, 70371, 70371, 70371, 70336, 70336, 70336, 70308, 70308, 70308, 70272, 70272, 70272, 70244, 70244, 70244, 70208, 70208, 70208, 70180, 70180, 70180, 70145, 70145, 70145, 70117, 70117, 70117, 70081, 70081, 70081, 70053, 70053, 70053, 70018, 70018, 70018, 69989, 69989, 69989, 69954, 69954, 69954, 69926, 69926, 69926, 69891, 69891, 69891, 69862, 69862, 69862, 69827, 69827, 69827, 69799, 69799, 69799, 69764, 69764, 69764, 69736, 69736, 69736, 69701, 69701, 69701, 69672, 69672, 69672, 69637, 69637, 69637, 69609, 69609, 69609, 69574, 69574, 69574, 69546, 69546, 69546, 69511, 69511, 69511, 69483, 69483, 69483, 69448, 69448, 69448, 69420, 69420, 69420, 69385, 69385, 69385, 69357, 69357, 69357, 69322, 69322, 69322, 69294, 69294, 69294, 69259, 69259, 69259, 69231, 69231, 69231, 69196, 69196, 69196, 69168, 69168, 69168, 69140, 69140, 69140, 69105, 69105, 69105, 69077, 69077, 69077, 69043, 69043, 69043, 69015, 69015, 69015, 68980, 68980, 68980, 68952, 68952, 68952, 68917, 68917, 68917, 68889, 68889, 68889, 68855, 68855, 68855, 68827, 68827, 68827, 68792, 68792, 68792, 68764, 68764, 68764, 68730, 68730, 68730, 68702, 68702, 68702, 68702, 68667, 68667, 68667, 68639, 68639, 68639, 68605, 68605, 68605, 68577, 68577, 68577, 68542, 68542, 68542, 68515, 68515, 68515, 68480, 68480, 68480, 68452, 68452, 68452, 68418, 68418, 68418, 68390, 68390, 68390, 68356, 68356, 68356, 68328, 68328, 68328, 68294, 68294, 68294, 68266, 68266, 68266, 68231, 68231, 68231, 68204, 68204, 68204, 68169, 68169, 68169, 68142, 68142, 68142, 68107, 68107, 68107, 68080, 68080, 68080, 68046, 68046, 68046, 68018, 68018, 68018, 67984, 67984, 67984, 67956, 67956, 67922, 67922, 67922, 67894, 67894, 67894, 67860, 67860, 67860, 67833, 67833, 67833, 67798, 67798, 67798, 67771, 67771, 67771, 67743, 67743, 67743, 67709, 67709, 67709, 67682, 67682, 67682, 67648, 67648, 67648, 67620, 67620, 67620, 67586, 67586, 67586, 67559, 67559, 67559, 67525, 67525, 67525, 67497, 67497, 67497, 67463, 67463, 67463, 67436, 67436, 67436, 67402, 67402, 67402, 67374, 67374, 67374, 67340, 67340, 67340, 67313, 67313, 67313, 67279, 67279, 67279, 67252, 67252, 67252, 67218, 67218, 67218, 67190, 67190, 67190, 67156, 67156, 67156, 67129, 67129, 67129, 67095, 67095, 67095, 67068, 67068, 67068, 67034, 67034, 67034, 67007, 67007, 67007, 66973, 66973, 66973, 66946, 66946, 66946, 66912, 66912, 66912, 66885, 66885, 66885, 66851, 66851, 66851, 66824, 66824, 66824, 66790, 66790, 66790, 66763, 66763, 66763, 66729, 66729, 66729, 66702, 66702, 66702, 66668, 66668, 66668, 66641, 66641, 66641, 66608, 66608, 66608, 66581, 66581, 66581, 66547, 66547, 66547, 66520, 66520, 66520, 66486, 66486, 66486, 66459, 66459, 66459, 66425, 66425, 66425, 66399, 66399, 66399, 66372, 66372, 66372, 66338, 66338, 66338, 66311, 66311, 66311, 66277, 66277, 66277, 66250, 66250, 66250, 66217, 66217, 66217, 66190, 66190, 66190, 66156, 66156, 66156, 66130, 66130, 66130, 66096, 66096, 66096, 66069, 66069, 66069, 66036, 66036, 66036, 66009, 66009, 66009, 65975, 65975, 65975, 65949, 65949, 65949, 65915, 65915, 65915, 65888, 65888, 65888, 65855, 65855, 65855, 65828, 65828, 65828, 65795, 65795, 65795, 65768, 65768, 65768, 65735, 65735, 65735, 65708, 65708, 65708, 65674, 65674, 65674, 65648, 65648, 65648, 65614, 65614, 65614, 65588, 65588, 65588, 65554, 65554, 65554, 65528, 65528, 65494, 65494, 65494, 65468, 65468, 65468, 65435, 65435, 65435, 65408, 65408, 65408, 65375, 65375, 65375, 65348, 65348, 65348, 65315, 65315, 65315, 65288, 65288, 65288, 65255, 65255, 65255, 65229, 65229, 65229, 65195, 65195, 65195, 65169, 65169, 65169, 65136, 65136, 65136, 65109, 65109, 65109, 65076, 65076, 65076, 65050, 65050, 65050, 65023, 65023, 65023, 64990, 64990, 64990, 64964, 64964, 64964, 64930, 64930, 64930, 64904, 64904, 64904, 64871, 64871, 64871, 64845, 64845, 64845, 64812, 64812, 64812, 64785, 64785, 64785, 64752, 64752, 64752, 64726, 64726, 64726, 64693, 64693, 64693, 64666, 64666, 64666, 64633, 64633, 64633, 64607, 64607, 64607, 64574, 64574, 64574, 64548, 64548, 64548, 64515, 64515, 64515, 64489, 64489, 64489, 64456, 64456, 64456, 64429, 64429, 64429, 64397, 64397, 64370, 64370, 64370, 64337, 64337, 64337, 64311, 64311, 64311, 64278, 64278, 64278, 64252, 64252, 64252, 64219, 64219, 64219, 64193, 64193, 64193, 64160, 64160, 64160, 64134, 64134, 64134, 64101, 64101, 64101, 64075, 64075, 64075, 64043, 64043, 64043, 64016, 64016, 64016, 63984, 63984, 63984, 63958, 63958, 63958, 63925, 63925, 63925, 63899, 63899, 63899, 63866, 63866, 63866, 63840, 63840, 63840, 63807, 63807, 63807, 63781, 63781, 63781, 63755, 63755, 63755, 63723, 63723, 63723, 63697, 63697, 63697, 63664, 63664, 63664, 63638, 63638, 63638, 63605, 63605, 63605, 63579, 63579, 63579, 63547, 63547, 63547, 63521, 63521, 63488, 63488, 63488, 63462, 63462, 63462, 63430, 63430, 63430, 63404, 63404, 63404, 63371, 63371, 63371, 63345, 63345, 63345, 63313, 63313, 63313, 63287, 63287, 63287, 63255, 63255, 63255, 63229, 63229, 63229, 63196, 63196, 63196, 63170, 63170, 63170, 63138, 63138, 63138, 63112, 63112, 63112, 63080, 63080, 63080, 63054, 63054, 63054, 63022, 63022, 63022, 62996, 62996, 62996, 62964, 62964, 62964, 62938, 62938, 62938, 62905, 62905, 62905, 62880, 62880, 62880, 62847, 62847, 62847, 62822, 62822, 62822, 62789, 62789, 62764, 62764, 62764, 62731, 62731, 62731, 62706, 62706, 62706, 62673, 62673, 62673, 62648, 62648, 62648, 62615, 62615, 62615, 62590, 62590, 62590, 62558, 62558, 62558, 62532, 62532, 62532, 62500, 62500, 62500, 62474, 62474, 62474, 62448, 62448, 62448, 62416, 62416, 62416, 62391, 62391, 62391, 62359, 62359, 62359, 62333, 62333, 62333, 62301, 62301, 62301, 62275, 62275, 62275, 62243, 62243, 62243, 62218, 62218, 62218, 62186, 62186, 62186, 62160, 62160, 62160, 62128, 62128, 62102, 62102, 62102, 62070, 62070, 62070, 62045, 62045, 62045, 62013, 62013, 62013, 61987, 61987, 61987, 61955, 61955, 61955, 61930, 61930, 61930, 61898, 61898, 61898, 61872, 61872, 61872, 61841, 61841, 61841, 61815, 61815, 61815, 61783, 61783, 61783, 61758, 61758, 61758, 61726, 61726, 61726, 61700, 61700, 61700, 61669, 61669, 61669, 61643, 61643, 61643, 61611, 61611, 61611, 61586, 61586, 61586, 61554, 61554, 61554, 61529, 61529, 61497, 61497, 61497, 61472, 61472, 61472, 61440, 61440, 61440, 61414, 61414, 61414, 61383, 61383, 61383, 61357, 61357, 61357, 61326, 61326, 61326, 61300, 61300, 61300, 61269, 61269, 61269, 61243, 61243, 61243, 61212, 61212, 61212, 61186, 61186, 61186, 61161, 61161, 61161, 61129, 61129, 61129, 61104, 61104, 61104, 61072, 61072, 61072, 61047, 61047, 61047, 61016, 61016, 61016, 60990, 60990, 60959, 60959, 60959, 60933, 60933, 60933, 60902, 60902, 60902, 60877, 60877, 60877, 60845, 60845, 60845, 60820, 60820, 60820, 60788, 60788, 60788, 60763, 60763, 60763, 60732, 60732, 60732, 60707, 60707, 60707, 60675, 60675, 60675, 60650, 60650, 60650, 60618, 60618, 60618, 60593, 60593, 60593, 60562, 60562, 60562, 60537, 60537, 60537, 60505, 60505, 60480, 60480, 60480, 60449, 60449, 60449, 60424, 60424, 60424, 60392, 60392, 60392, 60367, 60367, 60367, 60336, 60336, 60336, 60311, 60311, 60311, 60279, 60279, 60279, 60254, 60254, 60254, 60223, 60223, 60223, 60198, 60198, 60198, 60167, 60167, 60167, 60142, 60142, 60142, 60110, 60110, 60110, 60085, 60085, 60085, 60054, 60054, 60054, 60029, 60029, 59998, 59998, 59998, 59973, 59973, 59973, 59942, 59942, 59942, 59917, 59917, 59917, 59892, 59892, 59892, 59861, 59861, 59861, 59836, 59836, 59836, 59804, 59804, 59804, 59779, 59779, 59779, 59748, 59748, 59748, 59723, 59723, 59723, 59692, 59692, 59692, 59667, 59667, 59667, 59636, 59636, 59636, 59611, 59611, 59611, 59580, 59580, 59555, 59555, 59555, 59524, 59524, 59524, 59499, 59499, 59499, 59468, 59468, 59468, 59443, 59443, 59443, 59412, 59412, 59412, 59388, 59388, 59388, 59357, 59357, 59357, 59332, 59332, 59332, 59301, 59301, 59301, 59276, 59276, 59276, 59245, 59245, 59245, 59220, 59220, 59220, 59189, 59189, 59189, 59164, 59164, 59164, 59133, 59133, 59109, 59109, 59109, 59078, 59078, 59078, 59053, 59053, 59053, 59022, 59022, 59022, 58997, 58997, 58997, 58966, 58966, 58966, 58942, 58942, 58942, 58911, 58911, 58911, 58886, 58886, 58886, 58855, 58855, 58855, 58831, 58831, 58831, 58800, 58800, 58800, 58775, 58775, 58775, 58744, 58744, 58744, 58720, 58720, 58695, 58695, 58695, 58664, 58664, 58664, 58639, 58639, 58639, 58609, 58609, 58609, 58584, 58584, 58584, 58553, 58553, 58553, 58529, 58529, 58529, 58498, 58498, 58498, 58473, 58473, 58473, 58443, 58443, 58443, 58418, 58418, 58418, 58387, 58387, 58387, 58363, 58363, 58363, 58332, 58332, 58307, 58307, 58307, 58277, 58277, 58277, 58252, 58252, 58252, 58222, 58222, 58222, 58197, 58197, 58197, 58166, 58166, 58166, 58142, 58142, 58142, 58111, 58111, 58111, 58087, 58087, 58087, 58056, 58056, 58056, 58032, 58032, 58032, 58001, 58001, 58001, 57977, 57977, 57977, 57946, 57946, 57922, 57922, 57922, 57891, 57891, 57891, 57867, 57867, 57867, 57836, 57836, 57836, 57812, 57812, 57812, 57781, 57781, 57781, 57757, 57757, 57757, 57726, 57726, 57726, 57702, 57702, 57702, 57671, 57671, 57671, 57647, 57647, 57647, 57616, 57616, 57616, 57592, 57592, 57561, 57561, 57561, 57537, 57537, 57537, 57507, 57507, 57507, 57482, 57482, 57482, 57458, 57458, 57458, 57428, 57428, 57428, 57403, 57403, 57403, 57373, 57373, 57373, 57348, 57348, 57348, 57318, 57318, 57318, 57294, 57294, 57294, 57263, 57263, 57263, 57239, 57239, 57209, 57209, 57209, 57184, 57184, 57184, 57154, 57154, 57154, 57130, 57130, 57130, 57100, 57100, 57100, 57075, 57075, 57075, 57045, 57045, 57045, 57021, 57021, 57021, 56990, 56990, 56990, 56966, 56966, 56966, 56936, 56936, 56936, 56912, 56912, 56912, 56881, 56881, 56857, 56857, 56857, 56827, 56827, 56827, 56803, 56803, 56803, 56773, 56773, 56773, 56748, 56748, 56748, 56718, 56718, 56718, 56694, 56694, 56694, 56664, 56664, 56664, 56640, 56640, 56640, 56609, 56609, 56609, 56585, 56585, 56585, 56555, 56555, 56531, 56531, 56531, 56501, 56501, 56501, 56477, 56477, 56477, 56447, 56447, 56447, 56423, 56423, 56423, 56392, 56392, 56392, 56368, 56368, 56368, 56338, 56338, 56338, 56314, 56314, 56314, 56284, 56284, 56284, 56260, 56260, 56260, 56236, 56236, 56206, 56206, 56206, 56182, 56182, 56182, 56152, 56152, 56152, 56128, 56128, 56128, 56098, 56098, 56098, 56074, 56074, 56074, 56044, 56044, 56044, 56020, 56020, 56020, 55990, 55990, 55990, 55966, 55966, 55966, 55936, 55936, 55936, 55912, 55912, 55882, 55882, 55882, 55858, 55858, 55858, 55828, 55828, 55828, 55804, 55804, 55804, 55774, 55774, 55774, 55750, 55750, 55750, 55720, 55720, 55720, 55696, 55696, 55696, 55666, 55666, 55666, 55642, 55642, 55642, 55612, 55612, 55612, 55588, 55588, 55558, 55558, 55558, 55535, 55535, 55535, 55505, 55505, 55505, 55481, 55481, 55481, 55451, 55451, 55451, 55427, 55427, 55427, 55397, 55397, 55397, 55373, 55373, 55373, 55343, 55343, 55343, 55320, 55320, 55320, 55290, 55290, 55266, 55266, 55266, 55236, 55236, 55236, 55212, 55212, 55212, 55183, 55183, 55183, 55159, 55159, 55159, 55129, 55129, 55129, 55105, 55105, 55105, 55075, 55075, 55075, 55052, 55052, 55052, 55028, 55028, 55028, 54998, 54998, 54974, 54974, 54974, 54945, 54945, 54945, 54921, 54921, 54921, 54891, 54891, 54891, 54867, 54867, 54867, 54838, 54838, 54838, 54814, 54814, 54814, 54784, 54784, 54784, 54760, 54760, 54760, 54731, 54731, 54731, 54707, 54707, 54677, 54677, 54677, 54654, 54654, 54654, 54624, 54624, 54624, 54600, 54600, 54600, 54571, 54571, 54571, 54547, 54547, 54547, 54517, 54517, 54517, 54494, 54494, 54494, 54464, 54464, 54464, 54440, 54440, 54440, 54411, 54411, 54387, 54387, 54387, 54358, 54358, 54358, 54334, 54334, 54334, 54304, 54304, 54304, 54281, 54281, 54281, 54251, 54251, 54251, 54228, 54228, 54228, 54198, 54198, 54198, 54174, 54174, 54174, 54145, 54145, 54145, 54121, 54121, 54092, 54092, 54092, 54068, 54068, 54068, 54039, 54039, 54039, 54015, 54015, 54015, 53986, 53986, 53986, 53962, 53962, 53962, 53933, 53933, 53933, 53909, 53909, 53909, 53880, 53880, 53880, 53856, 53856, 53833, 53833, 53833, 53803, 53803, 53803, 53780, 53780, 53780, 53750, 53750, 53750, 53727, 53727, 53727, 53697, 53697, 53697, 53674, 53674, 53674, 53644, 53644, 53644, 53621, 53621, 53621, 53591, 53591, 53568, 53568, 53568, 53539, 53539, 53539, 53515, 53515, 53515, 53486, 53486, 53486, 53462, 53462, 53462, 53433, 53433, 53433, 53410, 53410, 53410, 53380, 53380, 53380, 53357, 53357, 53357, 53327, 53327, 53327, 53304, 53304, 53275, 53275, 53275, 53251, 53251, 53251, 53222, 53222, 53222, 53199, 53199, 53199, 53169, 53169, 53169, 53146, 53146, 53146, 53117, 53117, 53117, 53093, 53093, 53093, 53064, 53064, 53064, 53041, 53041, 53011, 53011, 53011, 52988, 52988, 52988, 52959, 52959, 52959, 52935, 52935, 52935, 52906, 52906, 52906, 52883, 52883, 52883, 52854, 52854, 52854, 52830, 52830, 52830, 52801, 52801, 52801, 52778, 52778, 52748, 52748, 52748, 52725, 52725, 52725, 52702, 52702, 52702, 52673, 52673, 52673, 52649, 52649, 52649, 52620, 52620, 52620, 52597, 52597, 52597, 52568, 52568, 52568, 52544, 52544, 52515, 52515, 52515, 52492, 52492, 52492, 52463, 52463, 52463, 52440, 52440, 52440, 52411, 52411, 52411, 52387, 52387, 52387, 52358, 52358, 52358, 52335, 52335, 52335, 52306, 52306, 52306, 52283, 52283, 52254, 52254, 52254, 52230, 52230, 52230, 52201, 52201, 52201, 52178, 52178, 52178, 52149, 52149, 52149, 52126, 52126, 52126, 52097, 52097, 52097, 52074, 52074, 52074, 52045, 52045, 52045, 52021, 52021, 51992, 51992, 51992, 51969, 51969, 51969, 51940, 51940, 51940, 51917, 51917, 51917, 51888, 51888, 51888, 51865, 51865, 51865, 51836, 51836, 51836, 51813, 51813, 51813, 51784, 51784, 51761, 51761, 51761, 51732, 51732, 51732, 51708, 51708, 51708, 51680, 51680, 51680, 51656, 51656, 51656, 51627, 51627, 51627, 51604, 51604, 51604, 51575, 51575, 51575, 51552, 51552, 51529, 51529, 51529, 51500, 51500, 51500, 51477, 51477, 51477, 51448, 51448, 51448, 51425, 51425, 51425, 51396, 51396, 51396, 51373, 51373, 51373, 51344, 51344, 51344, 51321, 51321, 51321, 51292, 51292, 51269, 51269, 51269, 51241, 51241, 51241, 51218, 51218, 51218, 51189, 51189, 51189, 51166, 51166, 51166, 51137, 51137, 51137, 51114, 51114, 51114, 51085, 51085, 51085, 51062, 51062, 51033, 51033, 51033, 51010, 51010, 51010, 50981, 50981, 50981, 50958, 50958, 50958, 50930, 50930, 50930, 50907, 50907, 50907, 50878, 50878, 50878, 50855, 50855, 50855, 50826, 50826, 50803, 50803, 50803, 50774, 50774, 50774, 50751, 50751, 50751, 50723, 50723, 50723, 50700, 50700, 50700, 50671, 50671, 50671, 50648, 50648, 50648, 50619, 50619, 50619, 50596, 50596, 50568, 50568, 50568, 50545, 50545, 50545, 50516, 50516, 50516, 50493, 50493, 50493, 50464, 50464, 50464, 50441, 50441, 50441, 50413, 50413, 50413, 50390, 50390, 50390, 50367, 50367, 50338, 50338, 50338, 50315, 50315, 50315, 50287, 50287, 50287, 50264, 50264, 50264, 50235, 50235, 50235, 50212, 50212, 50212, 50184, 50184, 50184, 50161, 50161, 50161, 50132, 50132, 50109, 50109, 50109, 50081, 50081, 50081, 50058, 50058, 50058, 50029, 50029, 50029, 50006, 50006, 50006, 49978, 49978, 49978, 49955, 49955, 49955, 49926, 49926, 49926, 49903, 49903, 49875, 49875, 49875, 49852, 49852, 49852, 49824, 49824, 49824, 49801, 49801, 49801, 49772, 49772, 49772, 49749, 49749, 49749, 49721, 49721, 49721, 49698, 49698, 49669, 49669, 49669, 49647, 49647, 49647, 49618, 49618, 49618, 49595, 49595, 49595, 49567, 49567, 49567, 49544, 49544, 49544, 49516, 49516, 49516, 49493, 49493, 49493, 49464, 49464, 49442, 49442, 49442, 49413, 49413, 49413, 49390, 49390, 49390, 49362, 49362, 49362, 49339, 49339, 49339, 49311, 49311, 49311, 49288, 49288, 49288, 49259, 49259, 49259, 49237, 49237, 49214, 49214, 49214, 49185, 49185, 49185, 49163, 49163, 49163, 49134, 49134, 49134, 49112, 49112, 49112, 49083, 49083, 49083, 49060, 49060, 49060, 49032, 49032, 49009, 49009, 49009, 48981, 48981, 48981, 48958, 48958, 48958, 48930, 48930, 48930, 48907, 48907, 48907, 48879, 48879, 48879, 48856, 48856, 48856, 48828, 48828, 48828, 48805, 48805, 48777, 48777, 48777, 48754, 48754, 48754, 48726, 48726, 48726, 48703, 48703, 48703, 48675, 48675, 48675, 48652, 48652, 48652, 48624, 48624, 48624, 48601, 48601, 48573, 48573, 48573, 48550, 48550, 48550, 48522, 48522, 48522, 48499, 48499, 48499, 48471, 48471, 48471, 48448, 48448, 48448, 48420, 48420, 48420, 48397, 48397, 48397, 48369, 48369, 48346, 48346, 48346, 48318, 48318, 48318, 48296, 48296, 48296, 48267, 48267, 48267, 48245, 48245, 48245, 48216, 48216, 48216, 48194, 48194, 48194, 48166, 48166, 48143, 48143, 48143, 48120, 48120, 48120, 48092, 48092, 48092, 48070, 48070, 48070, 48041, 48041, 48041, 48019, 48019, 48019, 47991, 47991, 47991, 47968, 47968, 47940, 47940, 47940, 47917, 47917, 47917, 47889, 47889, 47889, 47866, 47866, 47866, 47838, 47838, 47838, 47816, 47816, 47816, 47788, 47788, 47788, 47765, 47765, 47737, 47737, 47737, 47714, 47714, 47714, 47686, 47686, 47686, 47664, 47664, 47664, 47635, 47635, 47635, 47613, 47613, 47613, 47585, 47585, 47585, 47562, 47562, 47562, 47534, 47534, 47512, 47512, 47512, 47483, 47483, 47483, 47461, 47461, 47461, 47433, 47433, 47433, 47410, 47410, 47410, 47382, 47382, 47382, 47360, 47360, 47360, 47332, 47332, 47309, 47309, 47309, 47281, 47281, 47281, 47259, 47259, 47259, 47230, 47230, 47230, 47208, 47208, 47208, 47180, 47180, 47180, 47157, 47157, 47157, 47129, 47129, 47107, 47107, 47107, 47079, 47079, 47079, 47056, 47056, 47056, 47028, 47028, 47028, 47006, 47006, 47006, 46983, 46983, 46983, 46955, 46955, 46955, 46933, 46933, 46905, 46905, 46905, 46882, 46882, 46882, 46854, 46854, 46854, 46832, 46832, 46832, 46804, 46804, 46804, 46782, 46782, 46782, 46754, 46754, 46754, 46731, 46731, 46703, 46703, 46703, 46681, 46681, 46681, 46653, 46653, 46653, 46630, 46630, 46630, 46602, 46602, 46602, 46580, 46580, 46580, 46552, 46552, 46552, 46530, 46530, 46502, 46502, 46502, 46479, 46479, 46479, 46451, 46451, 46451, 46429, 46429, 46429, 46401, 46401, 46401, 46379, 46379, 46379, 46351, 46351, 46351, 46328, 46328, 46300, 46300, 46300, 46278, 46278, 46278, 46250, 46250, 46250, 46228, 46228, 46228, 46200, 46200, 46200, 46177, 46177, 46177, 46149, 46149, 46149, 46127, 46127, 46099, 46099, 46099, 46077, 46077, 46077, 46049, 46049, 46049, 46027, 46027, 46027, 45999, 45999, 45999, 45976, 45976, 45976, 45948, 45948, 45926, 45926, 45926, 45898, 45898, 45898, 45876, 45876, 45876, 45854, 45854, 45854, 45826, 45826, 45826, 45803, 45803, 45803, 45775, 45775, 45775, 45753, 45753, 45725, 45725, 45725, 45703, 45703, 45703, 45675, 45675, 45675, 45653, 45653, 45653, 45625, 45625, 45625, 45603, 45603, 45603, 45575, 45575, 45575, 45553, 45553, 45525, 45525, 45525, 45502, 45502, 45502, 45475, 45475, 45475, 45452, 45452, 45452, 45425, 45425, 45425, 45402, 45402, 45402, 45374, 45374, 45374, 45352, 45352, 45324, 45324, 45324, 45302, 45302, 45302, 45274, 45274, 45274, 45252, 45252, 45252, 45224, 45224, 45224, 45202, 45202, 45202, 45174, 45174, 45152, 45152, 45152, 45124, 45124, 45124, 45102, 45102, 45102, 45074, 45074, 45074, 45052, 45052, 45052, 45024, 45024, 45024, 45002, 45002, 45002, 44974, 44974, 44952, 44952, 44952, 44924, 44924, 44924, 44902, 44902, 44902, 44874, 44874, 44874, 44852, 44852, 44852, 44824, 44824, 44824, 44802, 44802, 44802, 44774, 44774, 44752, 44752, 44752, 44730, 44730, 44730, 44702, 44702, 44702, 44680, 44680, 44680, 44652, 44652, 44652, 44630, 44630, 44630, 44602, 44602, 44580, 44580, 44580, 44552, 44552, 44552, 44530, 44530, 44530, 44503, 44503, 44503, 44480, 44480, 44480, 44453, 44453, 44453, 44431, 44431, 44431, 44403, 44403, 44381, 44381, 44381, 44353, 44353, 44353, 44331, 44331, 44331, 44303, 44303, 44303, 44281, 44281, 44281, 44253, 44253, 44253, 44231, 44231, 44231, 44204, 44204, 44181, 44181, 44181, 44154, 44154, 44154, 44132, 44132, 44132, 44104, 44104, 44104, 44082, 44082, 44082, 44054, 44054, 44054, 44032, 44032, 44004, 44004, 44004, 43982, 43982, 43982, 43955, 43955, 43955, 43932, 43932, 43932, 43905, 43905, 43905, 43883, 43883, 43883, 43855, 43855, 43855, 43833, 43833, 43805, 43805, 43805, 43783, 43783, 43783, 43756, 43756, 43756, 43733, 43733, 43733, 43706, 43706, 43706, 43684, 43684, 43684, 43656, 43656, 43634, 43634, 43634, 43612, 43612, 43612, 43584, 43584, 43584, 43562, 43562, 43562, 43535, 43535, 43535, 43513, 43513, 43513, 43485, 43485, 43485, 43463, 43463, 43435, 43435, 43435, 43413, 43413, 43413, 43386, 43386, 43386, 43364, 43364, 43364, 43336, 43336, 43336, 43314, 43314, 43314, 43286, 43286, 43264, 43264, 43264, 43237, 43237, 43237, 43215, 43215, 43215, 43187, 43187, 43187, 43165, 43165, 43165, 43137, 43137, 43137, 43115, 43115, 43088, 43088, 43088, 43066, 43066, 43066, 43038, 43038, 43038, 43016, 43016, 43016, 42989, 42989, 42989, 42967, 42967, 42967, 42939, 42939, 42939, 42917, 42917, 42889, 42889, 42889, 42867, 42867, 42867, 42840, 42840, 42840, 42818, 42818, 42818, 42790, 42790, 42790, 42768, 42768, 42768, 42741, 42741, 42719, 42719, 42719, 42691, 42691, 42691, 42669, 42669, 42669, 42642, 42642, 42642, 42620, 42620, 42620, 42592, 42592, 42592, 42570, 42570, 42570, 42548, 42548, 42521, 42521, 42521, 42499, 42499, 42499, 42471, 42471, 42471, 42449, 42449, 42449, 42422, 42422, 42422, 42400, 42400, 42400, 42372, 42372, 42350, 42350, 42350, 42323, 42323, 42323, 42301, 42301, 42301, 42273, 42273, 42273, 42251, 42251, 42251, 42224, 42224, 42224, 42202, 42202, 42174, 42174, 42174, 42152, 42152, 42152, 42125, 42125, 42125, 42103, 42103, 42103, 42075, 42075, 42075, 42053, 42053, 42053, 42026, 42026, 42026, 42004, 42004, 41977, 41977, 41977, 41955, 41955, 41955, 41927, 41927, 41927, 41905, 41905, 41905, 41878, 41878, 41878, 41856, 41856, 41856, 41828, 41828, 41806, 41806, 41806, 41779, 41779, 41779, 41757, 41757, 41757, 41730, 41730, 41730, 41708, 41708, 41708, 41680, 41680, 41680, 41658, 41658, 41631, 41631, 41631, 41609, 41609, 41609, 41581, 41581, 41581, 41559, 41559, 41559, 41532, 41532, 41532, 41510, 41510, 41510, 41483, 41483, 41461, 41461, 41461, 41439, 41439, 41439, 41411, 41411, 41411, 41389, 41389, 41389, 41362, 41362, 41362, 41340, 41340, 41340, 41313, 41313, 41313, 41291, 41291, 41263, 41263, 41263, 41241, 41241, 41241, 41214, 41214, 41214, 41192, 41192, 41192, 41165, 41165, 41165, 41143, 41143, 41143, 41115, 41115, 41094, 41094, 41094, 41066, 41066, 41066, 41044, 41044, 41044, 41017, 41017, 41017, 40995, 40995, 40995, 40968, 40968, 40968, 40946, 40946, 40918, 40918, 40918, 40896, 40896, 40896, 40869, 40869, 40869, 40847, 40847, 40847, 40820, 40820, 40820, 40798, 40798, 40798, 40770, 40770, 40749, 40749, 40749, 40721, 40721, 40721, 40699, 40699, 40699, 40672, 40672, 40672, 40650, 40650, 40650, 40623, 40623, 40623, 40601, 40601, 40574, 40574, 40574, 40552, 40552, 40552, 40524, 40524, 40524, 40502, 40502, 40502, 40475, 40475, 40475, 40453, 40453, 40453, 40426, 40426, 40426, 40404, 40404, 40377, 40377, 40377, 40355, 40355, 40355, 40333, 40333, 40333, 40306, 40306, 40306, 40284, 40284, 40284, 40256, 40256, 40256, 40234, 40234, 40207, 40207, 40207, 40185, 40185, 40185, 40158, 40158, 40158, 40136, 40136, 40136, 40109, 40109, 40109, 40087, 40087, 40087, 40060, 40060, 40038, 40038, 40038, 40010, 40010, 40010, 39989, 39989, 39989, 39961, 39961, 39961, 39939, 39939, 39939, 39912, 39912, 39912, 39890, 39890, 39863, 39863, 39863, 39841, 39841, 39841, 39814, 39814, 39814, 39792, 39792, 39792, 39765, 39765, 39765, 39743, 39743, 39743, 39715, 39715, 39694, 39694, 39694, 39666, 39666, 39666, 39644, 39644, 39644, 39617, 39617, 39617, 39595, 39595, 39595, 39568, 39568, 39568, 39546, 39546, 39519, 39519, 39519, 39497, 39497, 39497, 39470, 39470, 39470, 39448, 39448, 39448, 39421, 39421, 39421, 39399, 39399, 39399, 39372, 39372, 39350, 39350, 39350, 39322, 39322, 39322, 39301, 39301, 39301, 39273, 39273, 39273, 39251, 39251, 39251, 39230, 39230, 39230, 39202, 39202, 39202, 39181, 39181, 39153, 39153, 39153, 39131, 39131, 39131, 39104, 39104, 39104, 39082, 39082, 39082, 39055, 39055, 39055, 39033, 39033, 39033, 39006, 39006, 38984, 38984, 38984, 38957, 38957, 38957, 38935, 38935, 38935, 38908, 38908, 38908, 38886, 38886, 38886, 38859, 38859, 38859, 38837, 38837, 38810, 38810, 38810, 38788, 38788, 38788, 38761, 38761, 38761, 38739, 38739, 38739, 38712, 38712, 38712, 38690, 38690, 38690, 38662, 38662, 38641, 38641, 38641, 38613, 38613, 38613, 38592, 38592, 38592, 38564, 38564, 38564, 38543, 38543, 38543, 38515, 38515, 38515, 38493, 38493, 38466, 38466, 38466, 38444, 38444, 38444, 38417, 38417, 38417, 38395, 38395, 38395, 38368, 38368, 38368, 38346, 38346, 38346, 38319, 38319, 38297, 38297, 38297, 38270, 38270, 38270, 38248, 38248, 38248, 38221, 38221, 38221, 38199, 38199, 38199, 38177, 38177, 38177, 38150, 38150, 38128, 38128, 38128, 38101, 38101, 38101, 38079, 38079, 38079, 38052, 38052, 38052, 38030, 38030, 38030, 38003, 38003, 38003, 37981, 37981, 37954, 37954, 37954, 37932, 37932, 37932, 37905, 37905, 37905, 37883, 37883, 37883, 37856, 37856, 37856, 37834, 37834, 37834, 37807, 37807, 37785, 37785, 37785, 37758, 37758, 37758, 37736, 37736, 37736, 37709, 37709, 37709, 37687, 37687, 37687, 37660, 37660, 37660, 37638, 37638, 37611, 37611, 37611, 37589, 37589, 37589, 37562, 37562, 37562, 37540, 37540, 37540, 37513, 37513, 37513, 37491, 37491, 37491, 37464, 37464, 37442, 37442, 37442, 37415, 37415, 37415, 37393, 37393, 37393, 37366, 37366, 37366, 37344, 37344, 37344, 37317, 37317, 37317, 37295, 37295, 37268, 37268, 37268, 37246, 37246, 37246, 37219, 37219, 37219, 37197, 37197, 37197, 37170, 37170, 37170, 37148, 37148, 37148, 37121, 37121, 37099, 37099, 37099, 37078, 37078, 37078, 37050, 37050, 37050, 37029, 37029, 37029, 37001, 37001, 37001, 36980, 36980, 36980, 36952, 36952, 36931, 36931, 36931, 36903, 36903, 36903, 36882, 36882, 36882, 36854, 36854, 36854, 36833, 36833, 36833, 36805, 36805, 36805, 36784, 36784, 36756, 36756, 36756, 36735, 36735, 36735, 36707, 36707, 36707, 36686, 36686, 36686, 36658, 36658, 36658, 36637, 36637, 36637, 36609, 36609, 36588, 36588, 36588, 36560, 36560, 36560, 36539, 36539, 36539, 36512, 36512, 36512, 36490, 36490, 36490, 36463, 36463, 36463, 36441, 36441, 36414, 36414, 36414, 36392, 36392, 36392, 36365, 36365, 36365, 36343, 36343, 36343, 36316, 36316, 36316, 36294, 36294, 36294, 36267, 36267, 36245, 36245, 36245, 36218, 36218, 36218, 36196, 36196, 36196, 36169, 36169, 36169, 36147, 36147, 36147, 36120, 36120, 36120, 36098, 36098, 36071, 36071, 36071, 36049, 36049, 36049, 36022, 36022, 36022, 36000, 36000);
    SIGNAL adc_sum_index : INTEGER RANGE 0 TO 72000;
BEGIN
    PROCESS (clk, rst)
    BEGIN
        IF rst = '1' THEN
            -- Reset the process if needed
            adc_sum_index <= 0;
        ELSIF rising_edge(clk) THEN
            -- Look up the adc_cum_sum in the LUT and get the corresponding index
            adc_sum_index <= lut_values(to_integer(adc_cum_sum));
        END IF;
    END PROCESS;

    -- Output the LUT index value
    lut_value <= adc_sum_index;
END main;